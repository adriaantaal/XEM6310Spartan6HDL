//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM, INC.
//Copyright (c) 2002-2011 ARM, Inc.
//The confidential and proprietary information contained in this file
//may only be used by a person authorised under and to the extent
//permitted by a subsisting licensing agreement from ARM Limited.
//
//(C) COPYRIGHT 2004-2011 ARM Limited.
//ALL RIGHTS RESERVED
//
//This entire notice must be reproduced on all copies of this file
//and copies of this file may only be made by a person if such person
//is permitted to do so under the terms of a subsisting license
//agreement from ARM Limited.
//

`ifdef ARM_UD_MODEL
`timescale 1ns/1ps
`define ARM_UD_DP  			#0.001
`define ARM_UD_DLY 			#0.02
`define ARM_UD_SEQ 			#0.01
`define ARM_UD_CP

`timescale 1ns/1ps
`celldefine
module ADDFHX1 (CO, S, A, B, CI);
output S, CO;
input A, B, CI;
  xor `ARM_UD_DP I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or `ARM_UD_DP I4(CO, a_and_b, a_and_ci, b_and_ci);
endmodule // ADDFHX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFHX2 (CO, S, A, B, CI);
output S, CO;
input A, B, CI;
  xor `ARM_UD_DP I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or `ARM_UD_DP I4(CO, a_and_b, a_and_ci, b_and_ci);
endmodule // ADDFHX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFHX4 (CO, S, A, B, CI);
output S, CO;
input A, B, CI;
  xor `ARM_UD_DP I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or `ARM_UD_DP I4(CO, a_and_b, a_and_ci, b_and_ci);
endmodule // ADDFHX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFHXL (CO, S, A, B, CI);
output S, CO;
input A, B, CI;
  xor `ARM_UD_DP I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or `ARM_UD_DP I4(CO, a_and_b, a_and_ci, b_and_ci);
endmodule // ADDFHXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFX1 (CO, S, A, B, CI);
output S, CO;
input A, B, CI;
  xor `ARM_UD_DP I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or `ARM_UD_DP I4(CO, a_and_b, a_and_ci, b_and_ci);
endmodule // ADDFX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFX2 (CO, S, A, B, CI);
output S, CO;
input A, B, CI;
  xor `ARM_UD_DP I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or `ARM_UD_DP I4(CO, a_and_b, a_and_ci, b_and_ci);
endmodule // ADDFX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFX4 (CO, S, A, B, CI);
output S, CO;
input A, B, CI;
  xor `ARM_UD_DP I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or `ARM_UD_DP I4(CO, a_and_b, a_and_ci, b_and_ci);
endmodule // ADDFX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFXL (CO, S, A, B, CI);
output S, CO;
input A, B, CI;
  xor `ARM_UD_DP I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or `ARM_UD_DP I4(CO, a_and_b, a_and_ci, b_and_ci);
endmodule // ADDFXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDHX1 (CO, S, A, B);
output S, CO;
input A, B;
  xor `ARM_UD_DP I0(S, A, B);
  and `ARM_UD_DP I1(CO, A, B);
endmodule // ADDHX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDHX2 (CO, S, A, B);
output S, CO;
input A, B;
  xor `ARM_UD_DP I0(S, A, B);
  and `ARM_UD_DP I1(CO, A, B);
endmodule // ADDHX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDHX4 (CO, S, A, B);
output S, CO;
input A, B;
  xor `ARM_UD_DP I0(S, A, B);
  and `ARM_UD_DP I1(CO, A, B);
endmodule // ADDHX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDHXL (CO, S, A, B);
output S, CO;
input A, B;
  xor `ARM_UD_DP I0(S, A, B);
  and `ARM_UD_DP I1(CO, A, B);
endmodule // ADDHXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AFCSHCINX2 (CO0, CO1, S, A, B, CI0N, CI1N, CS);
output S, CO0, CO1;
input A, B, CI0N, CI1N, CS;
  not I0 (cin1, CI1N);
  not I1 (cin0, CI0N);
  xor I2 (s1, A, B, cin1);
  xor I3 (s2, A, B, cin0);
  and I4 (s3, CS, s1);
  not I5 (csn, CS);
  and I6 (s4, csn, s2);
  or `ARM_UD_DP I7 (S, s3, s4);
  and I8 (a_and_b, A, B);
  and I9 (a_and_ci0, A, cin0);
  and I10 (b_and_ci0, B, cin0);
  or `ARM_UD_DP I11 (CO0, a_and_b, a_and_ci0, b_and_ci0);
  and I12 (a_and_ci1, A, cin1);
  and I13 (b_and_ci1, B, cin1);
  or `ARM_UD_DP I14 (CO1, a_and_b, a_and_ci1, b_and_ci1);
endmodule // AFCSHCINX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AFCSHCINX4 (CO0, CO1, S, A, B, CI0N, CI1N, CS);
output S, CO0, CO1;
input A, B, CI0N, CI1N, CS;
  not I0 (cin1, CI1N);
  not I1 (cin0, CI0N);
  xor I2 (s1, A, B, cin1);
  xor I3 (s2, A, B, cin0);
  and I4 (s3, CS, s1);
  not I5 (csn, CS);
  and I6 (s4, csn, s2);
  or `ARM_UD_DP I7 (S, s3, s4);
  and I8 (a_and_b, A, B);
  and I9 (a_and_ci0, A, cin0);
  and I10 (b_and_ci0, B, cin0);
  or `ARM_UD_DP I11 (CO0, a_and_b, a_and_ci0, b_and_ci0);
  and I12 (a_and_ci1, A, cin1);
  and I13 (b_and_ci1, B, cin1);
  or `ARM_UD_DP I14 (CO1, a_and_b, a_and_ci1, b_and_ci1);
endmodule // AFCSHCINX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AFCSHCONX2 (CO0N, CO1N, S, A, B, CI0, CI1, CS);
output S, CO0N, CO1N;
input A, B, CI0, CI1, CS;
  xor I2 (s1, A, B, CI1);
  xor I3 (s2, A, B, CI0);
  and I4 (s3, CS, s1);
  not I5 (csn, CS);
  and I6 (s4, csn, s2);
  or `ARM_UD_DP I7 (S, s3, s4);
  and I8 (a_and_b, A, B);
  and I9 (a_and_ci0, A, CI0);
  and I10 (b_and_ci0, B, CI0);
  or I11 (cout0, a_and_b, a_and_ci0, b_and_ci0);
  and I12 (a_and_ci1, A, CI1);
  and I13 (b_and_ci1, B, CI1);
  or I14 (cout1, a_and_b, a_and_ci1, b_and_ci1);
  not `ARM_UD_DP I15 (CO0N, cout0);
  not `ARM_UD_DP I16 (CO1N, cout1);
endmodule // AFCSHCONX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AFCSHCONX4 (CO0N, CO1N, S, A, B, CI0, CI1, CS);
output S, CO0N, CO1N;
input A, B, CI0, CI1, CS;
  xor I2 (s1, A, B, CI1);
  xor I3 (s2, A, B, CI0);
  and I4 (s3, CS, s1);
  not I5 (csn, CS);
  and I6 (s4, csn, s2);
  or `ARM_UD_DP I7 (S, s3, s4);
  and I8 (a_and_b, A, B);
  and I9 (a_and_ci0, A, CI0);
  and I10 (b_and_ci0, B, CI0);
  or I11 (cout0, a_and_b, a_and_ci0, b_and_ci0);
  and I12 (a_and_ci1, A, CI1);
  and I13 (b_and_ci1, B, CI1);
  or I14 (cout1, a_and_b, a_and_ci1, b_and_ci1);
  not `ARM_UD_DP I15 (CO0N, cout0);
  not `ARM_UD_DP I16 (CO1N, cout1);
endmodule // AFCSHCONX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AFHCINX2 (CO, S, A, B, CIN);
output S, CO;
input A, B, CIN;
  not I0 (ci, CIN);
  xor `ARM_UD_DP I1 (S, A, B, ci);
  and I2 (a_and_b, A, B);
  and I3 (a_and_ci, A, ci);
  and I4 (b_and_ci, B, ci);
  or `ARM_UD_DP I5 (CO, a_and_b, a_and_ci, b_and_ci);
endmodule // AFHCINX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AFHCINX4 (CO, S, A, B, CIN);
output S, CO;
input A, B, CIN;
  not I0 (ci, CIN);
  xor `ARM_UD_DP I1 (S, A, B, ci);
  and I2 (a_and_b, A, B);
  and I3 (a_and_ci, A, ci);
  and I4 (b_and_ci, B, ci);
  or `ARM_UD_DP I5 (CO, a_and_b, a_and_ci, b_and_ci);
endmodule // AFHCINX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AFHCONX2 (CON, S, A, B, CI);
output S, CON;
input A, B, CI;
  xor `ARM_UD_DP I0 (S, A, B, CI);
  and I1 (a_and_b, A, B);
  and I2 (a_and_ci, A, CI);
  and I3 (b_and_ci, B, CI);
  or I4 (cout, a_and_b, a_and_ci, b_and_ci);
  not `ARM_UD_DP I5 (CON, cout);
endmodule // AFHCONX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AFHCONX4 (CON, S, A, B, CI);
output S, CON;
input A, B, CI;
  xor `ARM_UD_DP I0 (S, A, B, CI);
  and I1 (a_and_b, A, B);
  and I2 (a_and_ci, A, CI);
  and I3 (b_and_ci, B, CI);
  or I4 (cout, a_and_b, a_and_ci, b_and_ci);
  not `ARM_UD_DP I5 (CON, cout);
endmodule // AFHCONX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AHHCINX2 (CO, S, A, CIN);
output S, CO;
input A, CIN;
  not I0 (ci, CIN);
  xor `ARM_UD_DP I1 (S, A, ci);
  and `ARM_UD_DP I2 (CO, A, ci);
endmodule // AHHCINX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AHHCINX4 (CO, S, A, CIN);
output S, CO;
input A, CIN;
  not I0 (ci, CIN);
  xor `ARM_UD_DP I1 (S, A, ci);
  and `ARM_UD_DP I2 (CO, A, ci);
endmodule // AHHCINX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AHHCONX2 (CON, S, A, CI);
output S, CON;
input A, CI;
  xor `ARM_UD_DP I0 (S, A, CI);
  and  I1 (cout, A, CI);
  not `ARM_UD_DP I2 (CON, cout);
endmodule // AHHCONX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AHHCONX4 (CON, S, A, CI);
output S, CON;
input A, CI;
  xor `ARM_UD_DP I0 (S, A, CI);
  and  I1 (cout, A, CI);
  not `ARM_UD_DP I2 (CON, cout);
endmodule // AHHCONX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2X1 (Y, A, B);
output Y;
input A, B;

  and `ARM_UD_DP (Y, A, B);
endmodule // AND2X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2X2 (Y, A, B);
output Y;
input A, B;

  and `ARM_UD_DP (Y, A, B);
endmodule // AND2X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2X4 (Y, A, B);
output Y;
input A, B;

  and `ARM_UD_DP (Y, A, B);
endmodule // AND2X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2XL (Y, A, B);
output Y;
input A, B;

  and `ARM_UD_DP (Y, A, B);
endmodule // AND2XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3X1 (Y, A, B, C);
output Y;
input A, B, C;

  and `ARM_UD_DP (Y, A, B, C);
endmodule // AND3X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3X2 (Y, A, B, C);
output Y;
input A, B, C;

  and `ARM_UD_DP (Y, A, B, C);
endmodule // AND3X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3X4 (Y, A, B, C);
output Y;
input A, B, C;

  and `ARM_UD_DP (Y, A, B, C);
endmodule // AND3X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3XL (Y, A, B, C);
output Y;
input A, B, C;

  and `ARM_UD_DP (Y, A, B, C);
endmodule // AND3XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4X1 (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and `ARM_UD_DP (Y, A, B, C, D);
endmodule // AND4X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4X2 (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and `ARM_UD_DP (Y, A, B, C, D);
endmodule // AND4X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4X4 (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and `ARM_UD_DP (Y, A, B, C, D);
endmodule // AND4X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4XL (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and `ARM_UD_DP (Y, A, B, C, D);
endmodule // AND4XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ANTENNA (A);
input A;
endmodule // ANTENNA
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211X1 (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor `ARM_UD_DP I1(Y, B0, C0, outA);
endmodule // AOI211X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211X2 (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor `ARM_UD_DP I1(Y, B0, C0, outA);
endmodule // AOI211X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211X4 (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor `ARM_UD_DP I1(Y, B0, C0, outA);
endmodule // AOI211X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211XL (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor `ARM_UD_DP I1(Y, B0, C0, outA);
endmodule // AOI211XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21X1 (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor `ARM_UD_DP I1(Y, B0, outA);
endmodule // AOI21X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21X2 (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor `ARM_UD_DP I1(Y, B0, outA);
endmodule // AOI21X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21X4 (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor `ARM_UD_DP I1(Y, B0, outA);
endmodule // AOI21X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21XL (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor `ARM_UD_DP I1(Y, B0, outA);
endmodule // AOI21XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221X1 (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, C0, outB, outA);
endmodule // AOI221X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221X2 (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, C0, outB, outA);
endmodule // AOI221X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221X4 (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, C0, outB, outA);
endmodule // AOI221X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221XL (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, C0, outB, outA);
endmodule // AOI221XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222X1 (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor `ARM_UD_DP I3(Y, outA, outB, outC);
endmodule // AOI222X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222X2 (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor `ARM_UD_DP I3(Y, outA, outB, outC);
endmodule // AOI222X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222X4 (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor `ARM_UD_DP I3(Y, outA, outB, outC);
endmodule // AOI222X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222XL (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor `ARM_UD_DP I3(Y, outA, outB, outC);
endmodule // AOI222XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22X1 (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, outA, outB);
endmodule // AOI22X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22X2 (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, outA, outB);
endmodule // AOI22X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22X4 (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, outA, outB);
endmodule // AOI22X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22XL (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, outA, outB);
endmodule // AOI22XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB1X1 (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;



  nor I0 (outA, A0N, A1N);
  nor `ARM_UD_DP I1 (Y, B0, outA);
endmodule // AOI2BB1X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB1X2 (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;



  nor I0 (outA, A0N, A1N);
  nor `ARM_UD_DP I1 (Y, B0, outA);
endmodule // AOI2BB1X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB1X4 (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;



  nor I0 (outA, A0N, A1N);
  nor `ARM_UD_DP I1 (Y, B0, outA);
endmodule // AOI2BB1X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB1XL (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;



  nor I0 (outA, A0N, A1N);
  nor `ARM_UD_DP I1 (Y, B0, outA);
endmodule // AOI2BB1XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB2X1 (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;



  nor I0 (outA, A0N, A1N);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, outA, outB);
endmodule // AOI2BB2X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB2X2 (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;



  nor I0 (outA, A0N, A1N);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, outA, outB);
endmodule // AOI2BB2X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB2X4 (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;



  nor I0 (outA, A0N, A1N);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, outA, outB);
endmodule // AOI2BB2X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB2XL (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;



  nor I0 (outA, A0N, A1N);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, outA, outB);
endmodule // AOI2BB2XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31X1 (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor `ARM_UD_DP I1(Y, B0, outA);
endmodule // AOI31X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31X2 (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor `ARM_UD_DP I1(Y, B0, outA);
endmodule // AOI31X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31X4 (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor `ARM_UD_DP I1(Y, B0, outA);
endmodule // AOI31X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31XL (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor `ARM_UD_DP I1(Y, B0, outA);
endmodule // AOI31XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32X1 (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, outA, outB);
endmodule // AOI32X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32X2 (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, outA, outB);
endmodule // AOI32X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32X4 (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, outA, outB);
endmodule // AOI32X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32XL (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor `ARM_UD_DP I2(Y, outA, outB);
endmodule // AOI32XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI33X1 (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1, B2);
  nor `ARM_UD_DP I2(Y, outA, outB);
endmodule // AOI33X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI33X2 (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1, B2);
  nor `ARM_UD_DP I2(Y, outA, outB);
endmodule // AOI33X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI33X4 (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1, B2);
  nor `ARM_UD_DP I2(Y, outA, outB);
endmodule // AOI33X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI33XL (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1, B2);
  nor `ARM_UD_DP I2(Y, outA, outB);
endmodule // AOI33XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BENCX1 (A, S, X2, M0, M1, M2);
output S, A, X2;
input M2, M1, M0;

  not I0 (m1n, M1);
  not I1 (m0n, M0);
  or  I3 (m1n_or_m0n, m1n, m0n);
  nand `ARM_UD_DP I4 (S, M2, m1n_or_m0n);
  or  I5 (m1_or_m0, M1, M0);
  nand `ARM_UD_DP I6 (A, m2n, m1_or_m0);
  xor I7 (x2n, M1, M0);
  not `ARM_UD_DP I8 (X2, x2n);
  not I9 (m2n, M2);

endmodule // BENCX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BENCX2 (A, S, X2, M0, M1, M2);
output S, A, X2;
input M2, M1, M0;

  not I0 (m1n, M1);
  not I1 (m0n, M0);
  or  I3 (m1n_or_m0n, m1n, m0n);
  nand `ARM_UD_DP I4 (S, M2, m1n_or_m0n);
  or  I5 (m1_or_m0, M1, M0);
  nand `ARM_UD_DP I6 (A, m2n, m1_or_m0);
  xor I7 (x2n, M1, M0);
  not `ARM_UD_DP I8 (X2, x2n);
  not I9 (m2n, M2);

endmodule // BENCX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BENCX4 (A, S, X2, M0, M1, M2);
output S, A, X2;
input M2, M1, M0;

  not I0 (m1n, M1);
  not I1 (m0n, M0);
  or  I3 (m1n_or_m0n, m1n, m0n);
  nand `ARM_UD_DP I4 (S, M2, m1n_or_m0n);
  or  I5 (m1_or_m0, M1, M0);
  nand `ARM_UD_DP I6 (A, m2n, m1_or_m0);
  xor I7 (x2n, M1, M0);
  not `ARM_UD_DP I8 (X2, x2n);
  not I9 (m2n, M2);

endmodule // BENCX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BMXX1 (PP, A, M0, M1, S, X2);
output PP;
input X2, A, S, M1, M0;

  udp_bmx `ARM_UD_DP I0 (PP, X2, A, S, M1, M0);

endmodule // BMXX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFX1 (Y, A);
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUFX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFX12 (Y, A);
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUFX12
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFX16 (Y, A);
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUFX16
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFX2 (Y, A);
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUFX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFX20 (Y, A);
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUFX20
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFX3 (Y, A);
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUFX3
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFX4 (Y, A);
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUFX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFX8 (Y, A);
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUFX8
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFXL (Y, A);
output Y;
input A;

  buf `ARM_UD_DP I0(Y, A);

endmodule // BUFXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUFX1 (Y, A);
output Y;
input A;

  buf `ARM_UD_CP I0(Y, A);

endmodule // CLKBUFX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUFX12 (Y, A);
output Y;
input A;

  buf `ARM_UD_CP I0(Y, A);

endmodule // CLKBUFX12
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUFX16 (Y, A);
output Y;
input A;

  buf `ARM_UD_CP I0(Y, A);

endmodule // CLKBUFX16
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUFX2 (Y, A);
output Y;
input A;

  buf `ARM_UD_CP I0(Y, A);

endmodule // CLKBUFX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUFX20 (Y, A);
output Y;
input A;

  buf `ARM_UD_CP I0(Y, A);

endmodule // CLKBUFX20
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUFX3 (Y, A);
output Y;
input A;

  buf `ARM_UD_CP I0(Y, A);

endmodule // CLKBUFX3
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUFX4 (Y, A);
output Y;
input A;

  buf `ARM_UD_CP I0(Y, A);

endmodule // CLKBUFX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUFX8 (Y, A);
output Y;
input A;

  buf `ARM_UD_CP I0(Y, A);

endmodule // CLKBUFX8
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUFXL (Y, A);
output Y;
input A;

  buf `ARM_UD_CP I0(Y, A);

endmodule // CLKBUFXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINVX1 (Y, A);
output Y;
input A;

  not `ARM_UD_CP I0(Y, A);

endmodule // CLKINVX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINVX12 (Y, A);
output Y;
input A;

  not `ARM_UD_CP I0(Y, A);

endmodule // CLKINVX12
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINVX16 (Y, A);
output Y;
input A;

  not `ARM_UD_CP I0(Y, A);

endmodule // CLKINVX16
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINVX2 (Y, A);
output Y;
input A;

  not `ARM_UD_CP I0(Y, A);

endmodule // CLKINVX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINVX20 (Y, A);
output Y;
input A;

  not `ARM_UD_CP I0(Y, A);

endmodule // CLKINVX20
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINVX3 (Y, A);
output Y;
input A;

  not `ARM_UD_CP I0(Y, A);

endmodule // CLKINVX3
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINVX4 (Y, A);
output Y;
input A;

  not `ARM_UD_CP I0(Y, A);

endmodule // CLKINVX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINVX8 (Y, A);
output Y;
input A;

  not `ARM_UD_CP I0(Y, A);

endmodule // CLKINVX8
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINVXL (Y, A);
output Y;
input A;

  not `ARM_UD_CP I0(Y, A);

endmodule // CLKINVXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CMPR22X1 (CO, S, A, B);
output S, CO;
input A, B;
  xor `ARM_UD_DP I0(S, A, B);
  and `ARM_UD_DP I1(CO, A, B);
endmodule // CMPR22X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CMPR32X1 (CO, S, A, B, C);
output S, CO;
input A, B, C;

  xor I0 (t1, A, B);
  xor `ARM_UD_DP I1 (S, t1, C);
  and I2 (t2, A, B);
  and I3 (t3, t1, C);
  or  `ARM_UD_DP I4 (CO, t2, t3);

endmodule // CMPR32X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CMPR42X1 (CO, ICO, S, A, B, C, D, ICI);
output S, CO, ICO;
input A, B, C, D, ICI;

  xor I0 (t1, A, B);
  xor I1 (IS, t1, C);
  and I2 (t2, A, B);
  and I3 (t3, A, C);
  and I4 (t4, B, C);
  or  `ARM_UD_DP  I5 (ICO, t2, t3, t4);
  xor I6 (ss, IS, D);
  xor `ARM_UD_DP  I7 (S, ss, ICI);
  and I8 (t5, IS, D);
  and I9 (t6, IS, ICI);
  and I10 (t7, D, ICI);
  or  `ARM_UD_DP  I11 (CO, t5, t6, t7);

endmodule // CMPR42X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CMPR42X2 (CO, ICO, S, A, B, C, D, ICI);
output S, CO, ICO;
input A, B, C, D, ICI;

  xor I0 (t1, A, B);
  xor I1 (IS, t1, C);
  and I2 (t2, A, B);
  and I3 (t3, A, C);
  and I4 (t4, B, C);
  or  `ARM_UD_DP  I5 (ICO, t2, t3, t4);
  xor I6 (ss, IS, D);
  xor `ARM_UD_DP  I7 (S, ss, ICI);
  and I8 (t5, IS, D);
  and I9 (t6, IS, ICI);
  and I10 (t7, D, ICI);
  or  `ARM_UD_DP  I11 (CO, t5, t6, t7);

endmodule // CMPR42X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DFFHQX1 (Q, CK, D);
output Q;
input  D, CK;
supply1 xSN,xRN;
  udp_dff_PWR I0 (n0, D, CK, xRN, xSN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFHQX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFHQX2 (Q, CK, D);
output Q;
input  D, CK;
supply1 xSN,xRN;
  udp_dff_PWR I0 (n0, D, CK, xRN, xSN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFHQX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFHQX4 (Q, CK, D);
output Q;
input  D, CK;
supply1 xSN,xRN;
  udp_dff_PWR I0 (n0, D, CK, xRN, xSN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFHQX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFHQXL (Q, CK, D);
output Q;
input  D, CK;
supply1 xSN,xRN;
  udp_dff_PWR I0 (n0, D, CK, xRN, xSN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFHQXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNRX1 (Q, QN, CKN, D, RN);
output Q, QN;
input  D, CKN, RN;
supply1 xSN;

  not      IC (clk, CKN);
  udp_dff_PWR I0 (n0, D, clk, RN, xSN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFNRX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNRX2 (Q, QN, CKN, D, RN);
output Q, QN;
input  D, CKN, RN;
supply1 xSN;

  not      IC (clk, CKN);
  udp_dff_PWR I0 (n0, D, clk, RN, xSN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFNRX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNRX4 (Q, QN, CKN, D, RN);
output Q, QN;
input  D, CKN, RN;
supply1 xSN;

  not      IC (clk, CKN);
  udp_dff_PWR I0 (n0, D, clk, RN, xSN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFNRX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNRXL (Q, QN, CKN, D, RN);
output Q, QN;
input  D, CKN, RN;
supply1 xSN;

  not      IC (clk, CKN);
  udp_dff_PWR I0 (n0, D, clk, RN, xSN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFNRXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSRX1 (Q, QN, CKN, D, RN, SN);
output Q, QN;
input  D, CKN, SN, RN;
  not      IC (clk, CKN);
  udp_dff_PWR I0 (n0, D, clk, RN, SN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFNSRX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSRX2 (Q, QN, CKN, D, RN, SN);
output Q, QN;
input  D, CKN, SN, RN;
  not      IC (clk, CKN);
  udp_dff_PWR I0 (n0, D, clk, RN, SN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFNSRX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSRX4 (Q, QN, CKN, D, RN, SN);
output Q, QN;
input  D, CKN, SN, RN;
  not      IC (clk, CKN);
  udp_dff_PWR I0 (n0, D, clk, RN, SN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFNSRX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSRXL (Q, QN, CKN, D, RN, SN);
output Q, QN;
input  D, CKN, SN, RN;
  not      IC (clk, CKN);
  udp_dff_PWR I0 (n0, D, clk, RN, SN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFNSRXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSX1 (Q, QN, CKN, D, SN);
output Q, QN;
input  D, CKN, SN;
supply1 xRN;

  not      IC (clk, CKN);
  udp_dff_PWR I0 (n0, D, clk, xRN, SN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFNSX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSX2 (Q, QN, CKN, D, SN);
output Q, QN;
input  D, CKN, SN;
supply1 xRN;

  not      IC (clk, CKN);
  udp_dff_PWR I0 (n0, D, clk, xRN, SN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFNSX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSX4 (Q, QN, CKN, D, SN);
output Q, QN;
input  D, CKN, SN;
supply1 xRN;

  not      IC (clk, CKN);
  udp_dff_PWR I0 (n0, D, clk, xRN, SN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFNSX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSXL (Q, QN, CKN, D, SN);
output Q, QN;
input  D, CKN, SN;
supply1 xRN;

  not      IC (clk, CKN);
  udp_dff_PWR I0 (n0, D, clk, xRN, SN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFNSXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNX1 (Q, QN, CKN, D);
output Q, QN;
input  D, CKN;
supply1 xSN,xRN;
  not      IC (clk, CKN);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFNX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNX2 (Q, QN, CKN, D);
output Q, QN;
input  D, CKN;
supply1 xSN,xRN;
  not      IC (clk, CKN);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFNX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNX4 (Q, QN, CKN, D);
output Q, QN;
input  D, CKN;
supply1 xSN,xRN;
  not      IC (clk, CKN);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFNX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNXL (Q, QN, CKN, D);
output Q, QN;
input  D, CKN;
supply1 xSN,xRN;
  not      IC (clk, CKN);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFNXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRHQX1 (Q, CK, D, RN);
output Q;
input  D, CK, RN;
supply1 xSN;

  udp_dff_PWR I0 (n0, D, CK, RN, xSN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFRHQX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRHQX2 (Q, CK, D, RN);
output Q;
input  D, CK, RN;
supply1 xSN;

  udp_dff_PWR I0 (n0, D, CK, RN, xSN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFRHQX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRHQX4 (Q, CK, D, RN);
output Q;
input  D, CK, RN;
supply1 xSN;

  udp_dff_PWR I0 (n0, D, CK, RN, xSN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFRHQX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRHQXL (Q, CK, D, RN);
output Q;
input  D, CK, RN;
supply1 xSN;

  udp_dff_PWR I0 (n0, D, CK, RN, xSN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFRHQXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRX1 (Q, QN, CK, D, RN);
output Q, QN;
input  D, CK, RN;
supply1 xSN;

  udp_dff_PWR I0 (n0, D, CK, RN, xSN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFRX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRX2 (Q, QN, CK, D, RN);
output Q, QN;
input  D, CK, RN;
supply1 xSN;

  udp_dff_PWR I0 (n0, D, CK, RN, xSN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFRX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRX4 (Q, QN, CK, D, RN);
output Q, QN;
input  D, CK, RN;
supply1 xSN;

  udp_dff_PWR I0 (n0, D, CK, RN, xSN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFRX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRXL (Q, QN, CK, D, RN);
output Q, QN;
input  D, CK, RN;
supply1 xSN;

  udp_dff_PWR I0 (n0, D, CK, RN, xSN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFRXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSHQX1 (Q, CK, D, SN);
output Q;
input  D, CK, SN;
supply1 xRN;

  udp_dff_PWR I0 (n0, D, CK, xRN, SN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFSHQX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSHQX2 (Q, CK, D, SN);
output Q;
input  D, CK, SN;
supply1 xRN;

  udp_dff_PWR I0 (n0, D, CK, xRN, SN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFSHQX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSHQX4 (Q, CK, D, SN);
output Q;
input  D, CK, SN;
supply1 xRN;

  udp_dff_PWR I0 (n0, D, CK, xRN, SN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFSHQX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSHQXL (Q, CK, D, SN);
output Q;
input  D, CK, SN;
supply1 xRN;

  udp_dff_PWR I0 (n0, D, CK, xRN, SN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFSHQXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRHQX1 (Q, CK, D, RN, SN);
output Q;
input  D, CK, SN, RN;
  udp_dff_PWR I0 (n0, D, CK, RN, SN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFSRHQX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRHQX2 (Q, CK, D, RN, SN);
output Q;
input  D, CK, SN, RN;
  udp_dff_PWR I0 (n0, D, CK, RN, SN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFSRHQX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRHQX4 (Q, CK, D, RN, SN);
output Q;
input  D, CK, SN, RN;
  udp_dff_PWR I0 (n0, D, CK, RN, SN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFSRHQX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRHQXL (Q, CK, D, RN, SN);
output Q;
input  D, CK, SN, RN;
  udp_dff_PWR I0 (n0, D, CK, RN, SN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
endmodule // DFFSRHQXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRX1 (Q, QN, CK, D, RN, SN);
output Q, QN;
input  D, CK, SN, RN;
  udp_dff_PWR I0 (n0, D, CK, RN, SN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFSRX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRX2 (Q, QN, CK, D, RN, SN);
output Q, QN;
input  D, CK, SN, RN;
  udp_dff_PWR I0 (n0, D, CK, RN, SN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFSRX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRX4 (Q, QN, CK, D, RN, SN);
output Q, QN;
input  D, CK, SN, RN;
  udp_dff_PWR I0 (n0, D, CK, RN, SN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFSRX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRXL (Q, QN, CK, D, RN, SN);
output Q, QN;
input  D, CK, SN, RN;
  udp_dff_PWR I0 (n0, D, CK, RN, SN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFSRXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSX1 (Q, QN, CK, D, SN);
output Q, QN;
input  D, CK, SN;
supply1 xRN;

  udp_dff_PWR I0 (n0, D, CK, xRN, SN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFSX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSX2 (Q, QN, CK, D, SN);
output Q, QN;
input  D, CK, SN;
supply1 xRN;

  udp_dff_PWR I0 (n0, D, CK, xRN, SN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFSX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSX4 (Q, QN, CK, D, SN);
output Q, QN;
input  D, CK, SN;
supply1 xRN;

  udp_dff_PWR I0 (n0, D, CK, xRN, SN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFSX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSXL (Q, QN, CK, D, SN);
output Q, QN;
input  D, CK, SN;
supply1 xRN;

  udp_dff_PWR I0 (n0, D, CK, xRN, SN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFSXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFTRX1 (Q, QN, CK, D, RN);
output Q, QN;
input  D, CK, RN;
supply1 xSN, EN,flag;

  udp_edfft_PWR I0 (n0, D, CK, RN, xSN, EN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFTRX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFTRX2 (Q, QN, CK, D, RN);
output Q, QN;
input  D, CK, RN;
supply1 xSN, EN,flag;

  udp_edfft_PWR I0 (n0, D, CK, RN, xSN, EN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFTRX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFTRX4 (Q, QN, CK, D, RN);
output Q, QN;
input  D, CK, RN;
supply1 xSN, EN,flag;

  udp_edfft_PWR I0 (n0, D, CK, RN, xSN, EN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFTRX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFTRXL (Q, QN, CK, D, RN);
output Q, QN;
input  D, CK, RN;
supply1 xSN, EN,flag;

  udp_edfft_PWR I0 (n0, D, CK, RN, xSN, EN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFTRXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFX1 (Q, QN, CK, D);
output Q, QN;
input  D, CK;
supply1 xSN,xRN;
  udp_dff_PWR I0 (n0, D, CK, xRN, xSN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFX2 (Q, QN, CK, D);
output Q, QN;
input  D, CK;
supply1 xSN,xRN;
  udp_dff_PWR I0 (n0, D, CK, xRN, xSN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFX4 (Q, QN, CK, D);
output Q, QN;
input  D, CK;
supply1 xSN,xRN;
  udp_dff_PWR I0 (n0, D, CK, xRN, xSN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFXL (Q, QN, CK, D);
output Q, QN;
input  D, CK;
supply1 xSN,xRN;
  udp_dff_PWR I0 (n0, D, CK, xRN, xSN, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // DFFXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DLY1X1 (Y, A);
output Y;
input A;

  buf `ARM_UD_DLY I0(Y, A);

endmodule // DLY1X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLY2X1 (Y, A);
output Y;
input A;

  buf `ARM_UD_DLY I0(Y, A);

endmodule // DLY2X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLY3X1 (Y, A);
output Y;
input A;

  buf `ARM_UD_DLY I0(Y, A);

endmodule // DLY3X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLY4X1 (Y, A);
output Y;
input A;

  buf `ARM_UD_DLY I0(Y, A);

endmodule // DLY4X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module EDFFTRX1 (Q, QN, CK, D, E, RN);
output Q, QN;
input D, CK, E, RN;
supply1 xSN;
supply1 dSN;

  udp_edfft_PWR I0 (n0, D, CK, RN, xSN, E, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // EDFFTRX1
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFFTRX2 (Q, QN, CK, D, E, RN);
output Q, QN;
input D, CK, E, RN;
supply1 xSN;
supply1 dSN;

  udp_edfft_PWR I0 (n0, D, CK, RN, xSN, E, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // EDFFTRX2
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFFTRX4 (Q, QN, CK, D, E, RN);
output Q, QN;
input D, CK, E, RN;
supply1 xSN;
supply1 dSN;

  udp_edfft_PWR I0 (n0, D, CK, RN, xSN, E, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // EDFFTRX4
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFFTRXL (Q, QN, CK, D, E, RN);
output Q, QN;
input D, CK, E, RN;
supply1 xSN;
supply1 dSN;

  udp_edfft_PWR I0 (n0, D, CK, RN, xSN, E, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ I1 (Q, n0);
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // EDFFTRXL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFFX1 (Q, QN, CK, D, E);
output Q, QN;
input D, CK, E;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff_PWR I0 (n0, D, CK, xRN, xSN, E, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ B1 (Q, n0);
  not      `ARM_UD_SEQ I1 (QN, n0);
endmodule // EDFFX1
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFFX2 (Q, QN, CK, D, E);
output Q, QN;
input D, CK, E;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff_PWR I0 (n0, D, CK, xRN, xSN, E, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ B1 (Q, n0);
  not      `ARM_UD_SEQ I1 (QN, n0);
endmodule // EDFFX2
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFFX4 (Q, QN, CK, D, E);
output Q, QN;
input D, CK, E;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff_PWR I0 (n0, D, CK, xRN, xSN, E, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ B1 (Q, n0);
  not      `ARM_UD_SEQ I1 (QN, n0);
endmodule // EDFFX4
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFFXL (Q, QN, CK, D, E);
output Q, QN;
input D, CK, E;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff_PWR I0 (n0, D, CK, xRN, xSN, E, 1'b1, 1'b0, 1'b1);
  buf     `ARM_UD_SEQ B1 (Q, n0);
  not      `ARM_UD_SEQ I1 (QN, n0);
endmodule // EDFFXL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module FILL1;
endmodule // FILL1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILL16;
endmodule // FILL16
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILL2;
endmodule // FILL2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILL32;
endmodule // FILL32
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILL4;
endmodule // FILL4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILL64;
endmodule // FILL64
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILL8;
endmodule // FILL8
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILLCAP16;
endmodule // FILLCAP16
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILLCAP3;
endmodule // FILLCAP3
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILLCAP32;
endmodule // FILLCAP32
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILLCAP4;
endmodule // FILLCAP4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILLCAP5;
endmodule // FILLCAP5
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILLCAP64;
endmodule // FILLCAP64
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILLCAP8;
endmodule // FILLCAP8
`endcelldefine
`timescale 1ns/1ps
`celldefine
module HOLDX1 (Y);
inout Y;

wire io_wire;

  buf(weak0,weak1) I0(Y, io_wire);
  buf I1(io_wire, Y);

endmodule // HOLDX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INVX1 (Y, A);
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INVX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INVX12 (Y, A);
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INVX12
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INVX16 (Y, A);
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INVX16
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INVX2 (Y, A);
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INVX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INVX20 (Y, A);
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INVX20
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INVX3 (Y, A);
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INVX3
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INVX4 (Y, A);
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INVX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INVX8 (Y, A);
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INVX8
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INVXL (Y, A);
output Y;
input A;

  not `ARM_UD_DP I0(Y, A);

endmodule // INVXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module JKFFRX1 (Q, QN, CK, J, K, RN);
output Q, QN;
input  J, K, CK, RN;
supply1 xSN;
supply1 dSN;


udp_jkff_PWR I0 (n0, J, K, CK, RN, xSN, 1'b1, 1'b0, 1'b1); 
buf `ARM_UD_SEQ I1 (Q,n0);
not `ARM_UD_SEQ I2 (QN,n0);

endmodule // JKFFRX1
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFRX2 (Q, QN, CK, J, K, RN);
output Q, QN;
input  J, K, CK, RN;
supply1 xSN;
supply1 dSN;


udp_jkff_PWR I0 (n0, J, K, CK, RN, xSN, 1'b1, 1'b0, 1'b1); 
buf `ARM_UD_SEQ I1 (Q,n0);
not `ARM_UD_SEQ I2 (QN,n0);

endmodule // JKFFRX2
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFRX4 (Q, QN, CK, J, K, RN);
output Q, QN;
input  J, K, CK, RN;
supply1 xSN;
supply1 dSN;


udp_jkff_PWR I0 (n0, J, K, CK, RN, xSN, 1'b1, 1'b0, 1'b1); 
buf `ARM_UD_SEQ I1 (Q,n0);
not `ARM_UD_SEQ I2 (QN,n0);

endmodule // JKFFRX4
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFRXL (Q, QN, CK, J, K, RN);
output Q, QN;
input  J, K, CK, RN;
supply1 xSN;
supply1 dSN;


udp_jkff_PWR I0 (n0, J, K, CK, RN, xSN, 1'b1, 1'b0, 1'b1); 
buf `ARM_UD_SEQ I1 (Q,n0);
not `ARM_UD_SEQ I2 (QN,n0);

endmodule // JKFFRXL
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFSRX1 (Q, QN, CK, J, K, RN, SN);
output Q, QN;
input  J, K, CK, SN, RN;


udp_jkff_PWR I0 (n0, J, K, CK, RN, SN, 1'b1, 1'b0, 1'b1); 
buf `ARM_UD_SEQ I1 (Q,n0);
not `ARM_UD_SEQ I2 (QN,n0);

endmodule // JKFFSRX1
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFSRX2 (Q, QN, CK, J, K, RN, SN);
output Q, QN;
input  J, K, CK, SN, RN;


udp_jkff_PWR I0 (n0, J, K, CK, RN, SN, 1'b1, 1'b0, 1'b1); 
buf `ARM_UD_SEQ I1 (Q,n0);
not `ARM_UD_SEQ I2 (QN,n0);

endmodule // JKFFSRX2
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFSRX4 (Q, QN, CK, J, K, RN, SN);
output Q, QN;
input  J, K, CK, SN, RN;


udp_jkff_PWR I0 (n0, J, K, CK, RN, SN, 1'b1, 1'b0, 1'b1); 
buf `ARM_UD_SEQ I1 (Q,n0);
not `ARM_UD_SEQ I2 (QN,n0);

endmodule // JKFFSRX4
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFSRXL (Q, QN, CK, J, K, RN, SN);
output Q, QN;
input  J, K, CK, SN, RN;


udp_jkff_PWR I0 (n0, J, K, CK, RN, SN, 1'b1, 1'b0, 1'b1); 
buf `ARM_UD_SEQ I1 (Q,n0);
not `ARM_UD_SEQ I2 (QN,n0);

endmodule // JKFFSRXL
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFSX1 (Q, QN, CK, J, K, SN);
output Q, QN;
input  J, K, CK, SN;
supply1 xRN;
supply1 dRN;

udp_jkff_PWR I0 (n0, J, K, CK, xRN, SN, 1'b1, 1'b0, 1'b1); 
buf `ARM_UD_SEQ I1 (Q,n0);
not `ARM_UD_SEQ I2 (QN,n0);

endmodule // JKFFSX1
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFSX2 (Q, QN, CK, J, K, SN);
output Q, QN;
input  J, K, CK, SN;
supply1 xRN;
supply1 dRN;

udp_jkff_PWR I0 (n0, J, K, CK, xRN, SN, 1'b1, 1'b0, 1'b1); 
buf `ARM_UD_SEQ I1 (Q,n0);
not `ARM_UD_SEQ I2 (QN,n0);

endmodule // JKFFSX2
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFSX4 (Q, QN, CK, J, K, SN);
output Q, QN;
input  J, K, CK, SN;
supply1 xRN;
supply1 dRN;

udp_jkff_PWR I0 (n0, J, K, CK, xRN, SN, 1'b1, 1'b0, 1'b1); 
buf `ARM_UD_SEQ I1 (Q,n0);
not `ARM_UD_SEQ I2 (QN,n0);

endmodule // JKFFSX4
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFSXL (Q, QN, CK, J, K, SN);
output Q, QN;
input  J, K, CK, SN;
supply1 xRN;
supply1 dRN;

udp_jkff_PWR I0 (n0, J, K, CK, xRN, SN, 1'b1, 1'b0, 1'b1); 
buf `ARM_UD_SEQ I1 (Q,n0);
not `ARM_UD_SEQ I2 (QN,n0);

endmodule // JKFFSXL
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFX1 (Q, QN, CK, J, K);
output Q, QN;
input  J, K, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;

udp_jkff_PWR I0 (n0, J, K, CK, xRN, xSN, 1'b1, 1'b0, 1'b1); 
buf `ARM_UD_SEQ I1 (Q,n0);
not `ARM_UD_SEQ I2 (QN,n0);

endmodule // JKFFX1
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFX2 (Q, QN, CK, J, K);
output Q, QN;
input  J, K, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;

udp_jkff_PWR I0 (n0, J, K, CK, xRN, xSN, 1'b1, 1'b0, 1'b1); 
buf `ARM_UD_SEQ I1 (Q,n0);
not `ARM_UD_SEQ I2 (QN,n0);

endmodule // JKFFX2
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFX4 (Q, QN, CK, J, K);
output Q, QN;
input  J, K, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;

udp_jkff_PWR I0 (n0, J, K, CK, xRN, xSN, 1'b1, 1'b0, 1'b1); 
buf `ARM_UD_SEQ I1 (Q,n0);
not `ARM_UD_SEQ I2 (QN,n0);

endmodule // JKFFX4
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFXL (Q, QN, CK, J, K);
output Q, QN;
input  J, K, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;

udp_jkff_PWR I0 (n0, J, K, CK, xRN, xSN, 1'b1, 1'b0, 1'b1); 
buf `ARM_UD_SEQ I1 (Q,n0);
not `ARM_UD_SEQ I2 (QN,n0);

endmodule // JKFFXL
`endcelldefine





`timescale 1ns/1ps
`celldefine
module MX2X1 (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MX2X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2X2 (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MX2X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2X4 (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MX2X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2XL (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 `ARM_UD_DP u0(Y, A, B, S0);

endmodule // MX2XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX4X1 (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 `ARM_UD_DP u0(Y, A, B, C, D, S0, S1);

endmodule // MX4X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX4X2 (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 `ARM_UD_DP u0(Y, A, B, C, D, S0, S1);

endmodule // MX4X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX4X4 (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 `ARM_UD_DP u0(Y, A, B, C, D, S0, S1);

endmodule // MX4X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX4XL (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 `ARM_UD_DP u0(Y, A, B, C, D, S0, S1);

endmodule // MX4XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2X1 (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      `ARM_UD_DP u1(Y, YN);

endmodule // MXI2X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2X2 (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      `ARM_UD_DP u1(Y, YN);

endmodule // MXI2X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2X4 (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      `ARM_UD_DP u1(Y, YN);

endmodule // MXI2X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2XL (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      `ARM_UD_DP u1(Y, YN);

endmodule // MXI2XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI4X1 (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      `ARM_UD_DP u1(Y, YN);

endmodule // MXI4X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI4X2 (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      `ARM_UD_DP u1(Y, YN);

endmodule // MXI4X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI4X4 (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      `ARM_UD_DP u1(Y, YN);

endmodule // MXI4X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI4XL (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      `ARM_UD_DP u1(Y, YN);

endmodule // MXI4XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2BX1 (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B);
endmodule // NAND2BX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2BX2 (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B);
endmodule // NAND2BX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2BX4 (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B);
endmodule // NAND2BX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2BXL (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B);
endmodule // NAND2BXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2X1 (Y, A, B);
output Y;
input A, B;

  nand `ARM_UD_DP (Y, A, B);
endmodule // NAND2X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2X2 (Y, A, B);
output Y;
input A, B;

  nand `ARM_UD_DP (Y, A, B);
endmodule // NAND2X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2X4 (Y, A, B);
output Y;
input A, B;

  nand `ARM_UD_DP (Y, A, B);
endmodule // NAND2X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2XL (Y, A, B);
output Y;
input A, B;

  nand `ARM_UD_DP (Y, A, B);
endmodule // NAND2XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BX1 (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B, C);
endmodule // NAND3BX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BX2 (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B, C);
endmodule // NAND3BX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BX4 (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B, C);
endmodule // NAND3BX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BXL (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B, C);
endmodule // NAND3BXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3X1 (Y, A, B, C);
output Y;
input A, B, C;

  nand `ARM_UD_DP (Y, A, B, C);
endmodule // NAND3X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3X2 (Y, A, B, C);
output Y;
input A, B, C;

  nand `ARM_UD_DP (Y, A, B, C);
endmodule // NAND3X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3X4 (Y, A, B, C);
output Y;
input A, B, C;

  nand `ARM_UD_DP (Y, A, B, C);
endmodule // NAND3X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3XL (Y, A, B, C);
output Y;
input A, B, C;

  nand `ARM_UD_DP (Y, A, B, C);
endmodule // NAND3XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BBX1 (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, Bx, C, D);
endmodule // NAND4BBX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BBX2 (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, Bx, C, D);
endmodule // NAND4BBX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BBX4 (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, Bx, C, D);
endmodule // NAND4BBX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BBXL (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, Bx, C, D);
endmodule // NAND4BBXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BX1 (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B, C, D);
endmodule // NAND4BX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BX2 (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B, C, D);
endmodule // NAND4BX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BX4 (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B, C, D);
endmodule // NAND4BX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BXL (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand `ARM_UD_DP (Y, Ax, B, C, D);
endmodule // NAND4BXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4X1 (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand `ARM_UD_DP (Y, A, B, C, D);
endmodule // NAND4X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4X2 (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand `ARM_UD_DP (Y, A, B, C, D);
endmodule // NAND4X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4X4 (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand `ARM_UD_DP (Y, A, B, C, D);
endmodule // NAND4X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4XL (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand `ARM_UD_DP (Y, A, B, C, D);
endmodule // NAND4XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2BX1 (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, B);
endmodule // NOR2BX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2BX2 (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, B);
endmodule // NOR2BX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2BX4 (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, B);
endmodule // NOR2BX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2BXL (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, B);
endmodule // NOR2BXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2X1 (Y, A, B);
output Y;
input A, B;

  nor `ARM_UD_DP (Y, A, B);
endmodule // NOR2X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2X2 (Y, A, B);
output Y;
input A, B;

  nor `ARM_UD_DP (Y, A, B);
endmodule // NOR2X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2X4 (Y, A, B);
output Y;
input A, B;

  nor `ARM_UD_DP (Y, A, B);
endmodule // NOR2X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2XL (Y, A, B);
output Y;
input A, B;

  nor `ARM_UD_DP (Y, A, B);
endmodule // NOR2XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BX1 (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, B, C);
endmodule // NOR3BX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BX2 (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, B, C);
endmodule // NOR3BX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BX4 (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, B, C);
endmodule // NOR3BX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BXL (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, B, C);
endmodule // NOR3BXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3X1 (Y, A, B, C);
output Y;
input A, B, C;

  nor `ARM_UD_DP (Y, A, B, C);
endmodule // NOR3X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3X2 (Y, A, B, C);
output Y;
input A, B, C;

  nor `ARM_UD_DP (Y, A, B, C);
endmodule // NOR3X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3X4 (Y, A, B, C);
output Y;
input A, B, C;

  nor `ARM_UD_DP (Y, A, B, C);
endmodule // NOR3X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3XL (Y, A, B, C);
output Y;
input A, B, C;

  nor `ARM_UD_DP (Y, A, B, C);
endmodule // NOR3XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BBX1 (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, Bx, C, D);
endmodule // NOR4BBX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BBX2 (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, Bx, C, D);
endmodule // NOR4BBX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BBX4 (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, Bx, C, D);
endmodule // NOR4BBX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BBXL (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, Bx, C, D);
endmodule // NOR4BBXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BX1 (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, B, C, D);
endmodule // NOR4BX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BX2 (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, B, C, D);
endmodule // NOR4BX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BX4 (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, B, C, D);
endmodule // NOR4BX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BXL (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nor `ARM_UD_DP (Y, Ax, B, C, D);
endmodule // NOR4BXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4X1 (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nor `ARM_UD_DP (Y, A, B, C, D);
endmodule // NOR4X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4X2 (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nor `ARM_UD_DP (Y, A, B, C, D);
endmodule // NOR4X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4X4 (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nor `ARM_UD_DP (Y, A, B, C, D);
endmodule // NOR4X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4XL (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nor `ARM_UD_DP (Y, A, B, C, D);
endmodule // NOR4XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211X1 (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand `ARM_UD_DP I1(Y, B0, C0, outA);
endmodule // OAI211X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211X2 (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand `ARM_UD_DP I1(Y, B0, C0, outA);
endmodule // OAI211X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211X4 (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand `ARM_UD_DP I1(Y, B0, C0, outA);
endmodule // OAI211X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211XL (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand `ARM_UD_DP I1(Y, B0, C0, outA);
endmodule // OAI211XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21X1 (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand `ARM_UD_DP I1(Y, B0, outA);
endmodule // OAI21X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21X2 (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand `ARM_UD_DP I1(Y, B0, outA);
endmodule // OAI21X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21X4 (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand `ARM_UD_DP I1(Y, B0, outA);
endmodule // OAI21X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21XL (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand `ARM_UD_DP I1(Y, B0, outA);
endmodule // OAI21XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221X1 (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand `ARM_UD_DP I2(Y, C0, outB, outA);
endmodule // OAI221X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221X2 (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand `ARM_UD_DP I2(Y, C0, outB, outA);
endmodule // OAI221X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221X4 (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand `ARM_UD_DP I2(Y, C0, outB, outA);
endmodule // OAI221X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221XL (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand `ARM_UD_DP I2(Y, C0, outB, outA);
endmodule // OAI221XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222X1 (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand `ARM_UD_DP I3(Y, outA, outB, outC);
endmodule // OAI222X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222X2 (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand `ARM_UD_DP I3(Y, outA, outB, outC);
endmodule // OAI222X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222X4 (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand `ARM_UD_DP I3(Y, outA, outB, outC);
endmodule // OAI222X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222XL (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand `ARM_UD_DP I3(Y, outA, outB, outC);
endmodule // OAI222XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22X1 (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand `ARM_UD_DP I2(Y, outA, outB);
endmodule // OAI22X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22X2 (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand `ARM_UD_DP I2(Y, outA, outB);
endmodule // OAI22X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22X4 (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand `ARM_UD_DP I2(Y, outA, outB);
endmodule // OAI22X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22XL (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand `ARM_UD_DP I2(Y, outA, outB);
endmodule // OAI22XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB1X1 (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;



  nand I0 (outA, A0N, A1N);
  nand `ARM_UD_DP I1(Y, B0, outA);
endmodule // OAI2BB1X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB1X2 (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;



  nand I0 (outA, A0N, A1N);
  nand `ARM_UD_DP I1(Y, B0, outA);
endmodule // OAI2BB1X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB1X4 (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;



  nand I0 (outA, A0N, A1N);
  nand `ARM_UD_DP I1(Y, B0, outA);
endmodule // OAI2BB1X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB1XL (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;



  nand I0 (outA, A0N, A1N);
  nand `ARM_UD_DP I1(Y, B0, outA);
endmodule // OAI2BB1XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB2X1 (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;



  nand I0 (outA, A0N, A1N);
  or   I1(outB, B0, B1);
  nand `ARM_UD_DP I2(Y, outA, outB);
endmodule // OAI2BB2X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB2X2 (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;



  nand I0 (outA, A0N, A1N);
  or   I1(outB, B0, B1);
  nand `ARM_UD_DP I2(Y, outA, outB);
endmodule // OAI2BB2X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB2X4 (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;



  nand I0 (outA, A0N, A1N);
  or   I1(outB, B0, B1);
  nand `ARM_UD_DP I2(Y, outA, outB);
endmodule // OAI2BB2X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB2XL (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;



  nand I0 (outA, A0N, A1N);
  or   I1(outB, B0, B1);
  nand `ARM_UD_DP I2(Y, outA, outB);
endmodule // OAI2BB2XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31X1 (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand `ARM_UD_DP I1(Y, B0, outA);
endmodule // OAI31X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31X2 (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand `ARM_UD_DP I1(Y, B0, outA);
endmodule // OAI31X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31X4 (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand `ARM_UD_DP I1(Y, B0, outA);
endmodule // OAI31X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31XL (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand `ARM_UD_DP I1(Y, B0, outA);
endmodule // OAI31XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI32X1 (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1);
  nand `ARM_UD_DP I2(Y, outA, outB);
endmodule // OAI32X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI32X2 (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1);
  nand `ARM_UD_DP I2(Y, outA, outB);
endmodule // OAI32X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI32X4 (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1);
  nand `ARM_UD_DP I2(Y, outA, outB);
endmodule // OAI32X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI32XL (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1);
  nand `ARM_UD_DP I2(Y, outA, outB);
endmodule // OAI32XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI33X1 (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1, B2);
  nand `ARM_UD_DP I2(Y, outA, outB);
endmodule // OAI33X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI33X2 (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1, B2);
  nand `ARM_UD_DP I2(Y, outA, outB);
endmodule // OAI33X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI33X4 (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1, B2);
  nand `ARM_UD_DP I2(Y, outA, outB);
endmodule // OAI33X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI33XL (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1, B2);
  nand `ARM_UD_DP I2(Y, outA, outB);
endmodule // OAI33XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2X1 (Y, A, B);
output Y;
input A, B;

  or `ARM_UD_DP (Y, A, B);
endmodule // OR2X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2X2 (Y, A, B);
output Y;
input A, B;

  or `ARM_UD_DP (Y, A, B);
endmodule // OR2X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2X4 (Y, A, B);
output Y;
input A, B;

  or `ARM_UD_DP (Y, A, B);
endmodule // OR2X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2XL (Y, A, B);
output Y;
input A, B;

  or `ARM_UD_DP (Y, A, B);
endmodule // OR2XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3X1 (Y, A, B, C);
output Y;
input A, B, C;

  or `ARM_UD_DP (Y, A, B, C);
endmodule // OR3X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3X2 (Y, A, B, C);
output Y;
input A, B, C;

  or `ARM_UD_DP (Y, A, B, C);
endmodule // OR3X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3X4 (Y, A, B, C);
output Y;
input A, B, C;

  or `ARM_UD_DP (Y, A, B, C);
endmodule // OR3X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3XL (Y, A, B, C);
output Y;
input A, B, C;

  or `ARM_UD_DP (Y, A, B, C);
endmodule // OR3XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4X1 (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or `ARM_UD_DP (Y, A, B, C, D);
endmodule // OR4X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4X2 (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or `ARM_UD_DP (Y, A, B, C, D);
endmodule // OR4X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4X4 (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or `ARM_UD_DP (Y, A, B, C, D);
endmodule // OR4X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4XL (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or `ARM_UD_DP (Y, A, B, C, D);
endmodule // OR4XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF1R1WX2 (RB, RW, RWN, WB, WW);
output RB;
input WB, WW, RW, RWN;

   not II (wwn,WW);
   udp_tlatrf I0 (n0, WB, WW, wwn, 1'b1);
   notif1     `ARM_UD_SEQ I1 (RB, n0, n2);
   udp_outrf  I2 (n2, n0, RWN, RW);




endmodule // RF1R1WX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF2R1WX2 (R1B, R2B, R1W, R2W, WB, WW);
output R1B, R2B;
input WB, WW, R1W, R2W;

   not        I0 (WWN, WW);
   not        I1 (R1WN, R1W);
   not        I2 (R2WN, R2W);
   udp_tlatrf I3 (n0, WB, WW, WWN, 1'b1);
   notif1     `ARM_UD_SEQ I4 (R1B, n0, n2);
   notif1     `ARM_UD_SEQ I5 (R2B, n0, n3);
   udp_outrf  I6 (n2, n0, R1WN, R1W);
   udp_outrf  I7 (n3, n0, R2WN, R2W);




endmodule // RF2R1WX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RFRDX1 (BRB, RB);
output BRB;
input RB;

   not(weak0,weak1) I0(RB, io_wire);
   not              I1(io_wire, RB);
   buf              `ARM_UD_SEQ I2(BRB, io_wire);




endmodule // RFRDX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RFRDX2 (BRB, RB);
output BRB;
input RB;

   not(weak0,weak1) I0(RB, io_wire);
   not              I1(io_wire, RB);
   buf              `ARM_UD_SEQ I2(BRB, io_wire);




endmodule // RFRDX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RFRDX4 (BRB, RB);
output BRB;
input RB;

   not(weak0,weak1) I0(RB, io_wire);
   not              I1(io_wire, RB);
   buf              `ARM_UD_SEQ I2(BRB, io_wire);




endmodule // RFRDX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RSLATNX1 (Q, QN, RN, SN);
output Q, QN;
input RN, SN;
  not I4(R, RN);
  not I5(S, SN);
  udp_rslat_pwr  I0(q,  R, S, 1'b1, 1'b0, 1'b1);
  udp_rslatn_pwr I1(qn, R, S, 1'b1, 1'b0, 1'b1);
  not `ARM_UD_SEQ I2(QN, q);
  not `ARM_UD_SEQ I3(Q, qn);

endmodule // RSLATNX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RSLATNX2 (Q, QN, RN, SN);
output Q, QN;
input RN, SN;
  not I4(R, RN);
  not I5(S, SN);
  udp_rslat_pwr  I0(q,  R, S, 1'b1, 1'b0, 1'b1);
  udp_rslatn_pwr I1(qn, R, S, 1'b1, 1'b0, 1'b1);
  not `ARM_UD_SEQ I2(QN, q);
  not `ARM_UD_SEQ I3(Q, qn);

endmodule // RSLATNX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RSLATNX4 (Q, QN, RN, SN);
output Q, QN;
input RN, SN;
  not I4(R, RN);
  not I5(S, SN);
  udp_rslat_pwr  I0(q,  R, S, 1'b1, 1'b0, 1'b1);
  udp_rslatn_pwr I1(qn, R, S, 1'b1, 1'b0, 1'b1);
  not `ARM_UD_SEQ I2(QN, q);
  not `ARM_UD_SEQ I3(Q, qn);

endmodule // RSLATNX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RSLATNXL (Q, QN, RN, SN);
output Q, QN;
input RN, SN;
  not I4(R, RN);
  not I5(S, SN);
  udp_rslat_pwr  I0(q,  R, S, 1'b1, 1'b0, 1'b1);
  udp_rslatn_pwr I1(qn, R, S, 1'b1, 1'b0, 1'b1);
  not `ARM_UD_SEQ I2(QN, q);
  not `ARM_UD_SEQ I3(Q, qn);

endmodule // RSLATNXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RSLATX1 (Q, QN, R, S);
output Q, QN;
input R, S;
  udp_rslat_pwr I0(q, R, S, 1'b1, 1'b0, 1'b1);
  udp_rslatn_pwr  I1(qn, R, S, 1'b1, 1'b0, 1'b1);
  buf `ARM_UD_SEQ I2(QN, qn);
  buf `ARM_UD_SEQ I3(Q, q);

endmodule // RSLATX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RSLATX2 (Q, QN, R, S);
output Q, QN;
input R, S;
  udp_rslat_pwr I0(q, R, S, 1'b1, 1'b0, 1'b1);
  udp_rslatn_pwr  I1(qn, R, S, 1'b1, 1'b0, 1'b1);
  buf `ARM_UD_SEQ I2(QN, qn);
  buf `ARM_UD_SEQ I3(Q, q);

endmodule // RSLATX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RSLATX4 (Q, QN, R, S);
output Q, QN;
input R, S;
  udp_rslat_pwr I0(q, R, S, 1'b1, 1'b0, 1'b1);
  udp_rslatn_pwr  I1(qn, R, S, 1'b1, 1'b0, 1'b1);
  buf `ARM_UD_SEQ I2(QN, qn);
  buf `ARM_UD_SEQ I3(Q, q);

endmodule // RSLATX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RSLATXL (Q, QN, R, S);
output Q, QN;
input R, S;
  udp_rslat_pwr I0(q, R, S, 1'b1, 1'b0, 1'b1);
  udp_rslatn_pwr  I1(qn, R, S, 1'b1, 1'b0, 1'b1);
  buf `ARM_UD_SEQ I2(QN, qn);
  buf `ARM_UD_SEQ I3(Q, q);

endmodule // RSLATXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module SDFFHQX1 (Q, CK, D, SE, SI);
output Q;
input D, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  udp_dff_PWR I0 (n0, n1, CK, xRN, xSN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFHQX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFHQX2 (Q, CK, D, SE, SI);
output Q;
input D, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  udp_dff_PWR I0 (n0, n1, CK, xRN, xSN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFHQX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFHQX4 (Q, CK, D, SE, SI);
output Q;
input D, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  udp_dff_PWR I0 (n0, n1, CK, xRN, xSN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFHQX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFHQXL (Q, CK, D, SE, SI);
output Q;
input D, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  udp_dff_PWR I0 (n0, n1, CK, xRN, xSN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFHQXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNRX1 (Q, QN, CKN, D, RN, SE, SI);
output Q, QN;
input D, SI, SE, CKN, RN;
supply1 xSN;
supply1 dSN;

  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, n1, clk, RN, xSN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFNRX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNRX2 (Q, QN, CKN, D, RN, SE, SI);
output Q, QN;
input D, SI, SE, CKN, RN;
supply1 xSN;
supply1 dSN;

  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, n1, clk, RN, xSN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFNRX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNRX4 (Q, QN, CKN, D, RN, SE, SI);
output Q, QN;
input D, SI, SE, CKN, RN;
supply1 xSN;
supply1 dSN;

  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, n1, clk, RN, xSN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFNRX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNRXL (Q, QN, CKN, D, RN, SE, SI);
output Q, QN;
input D, SI, SE, CKN, RN;
supply1 xSN;
supply1 dSN;

  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, n1, clk, RN, xSN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFNRXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSRX1 (Q, QN, CKN, D, RN, SE, SI, SN);
output Q, QN;
input D, SI, SE, CKN, SN, RN;
  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, n1, clk, RN, SN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFNSRX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSRX2 (Q, QN, CKN, D, RN, SE, SI, SN);
output Q, QN;
input D, SI, SE, CKN, SN, RN;
  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, n1, clk, RN, SN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFNSRX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSRX4 (Q, QN, CKN, D, RN, SE, SI, SN);
output Q, QN;
input D, SI, SE, CKN, SN, RN;
  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, n1, clk, RN, SN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFNSRX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSRXL (Q, QN, CKN, D, RN, SE, SI, SN);
output Q, QN;
input D, SI, SE, CKN, SN, RN;
  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, n1, clk, RN, SN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFNSRXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSX1 (Q, QN, CKN, D, SE, SI, SN);
output Q, QN;
input D, SI, SE, CKN, SN;
supply1 xRN;
supply1 dRN;

  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, n1, clk, xRN, SN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFNSX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSX2 (Q, QN, CKN, D, SE, SI, SN);
output Q, QN;
input D, SI, SE, CKN, SN;
supply1 xRN;
supply1 dRN;

  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, n1, clk, xRN, SN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFNSX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSX4 (Q, QN, CKN, D, SE, SI, SN);
output Q, QN;
input D, SI, SE, CKN, SN;
supply1 xRN;
supply1 dRN;

  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, n1, clk, xRN, SN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFNSX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSXL (Q, QN, CKN, D, SE, SI, SN);
output Q, QN;
input D, SI, SE, CKN, SN;
supply1 xRN;
supply1 dRN;

  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, n1, clk, xRN, SN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFNSXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNX1 (Q, QN, CKN, D, SE, SI);
output Q, QN;
input D, SI, SE, CKN;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFNX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNX2 (Q, QN, CKN, D, SE, SI);
output Q, QN;
input D, SI, SE, CKN;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFNX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNX4 (Q, QN, CKN, D, SE, SI);
output Q, QN;
input D, SI, SE, CKN;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFNX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNXL (Q, QN, CKN, D, SE, SI);
output Q, QN;
input D, SI, SE, CKN;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFNXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRHQX1 (Q, CK, D, RN, SE, SI);
output Q;
input D, SI, SE, CK, RN;
supply1 xSN;
supply1 dSN;

  udp_dff_PWR I0 (n0, n1, CK, RN, xSN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFRHQX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRHQX2 (Q, CK, D, RN, SE, SI);
output Q;
input D, SI, SE, CK, RN;
supply1 xSN;
supply1 dSN;

  udp_dff_PWR I0 (n0, n1, CK, RN, xSN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFRHQX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRHQX4 (Q, CK, D, RN, SE, SI);
output Q;
input D, SI, SE, CK, RN;
supply1 xSN;
supply1 dSN;

  udp_dff_PWR I0 (n0, n1, CK, RN, xSN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFRHQX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRHQXL (Q, CK, D, RN, SE, SI);
output Q;
input D, SI, SE, CK, RN;
supply1 xSN;
supply1 dSN;

  udp_dff_PWR I0 (n0, n1, CK, RN, xSN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFRHQXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRX1 (Q, QN, CK, D, RN, SE, SI);
output Q, QN;
input D, SI, SE, CK, RN;
supply1 xSN;
supply1 dSN;

  udp_dff_PWR I0 (n0, n1, CK, RN, xSN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFRX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRX2 (Q, QN, CK, D, RN, SE, SI);
output Q, QN;
input D, SI, SE, CK, RN;
supply1 xSN;
supply1 dSN;

  udp_dff_PWR I0 (n0, n1, CK, RN, xSN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFRX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRX4 (Q, QN, CK, D, RN, SE, SI);
output Q, QN;
input D, SI, SE, CK, RN;
supply1 xSN;
supply1 dSN;

  udp_dff_PWR I0 (n0, n1, CK, RN, xSN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFRX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRXL (Q, QN, CK, D, RN, SE, SI);
output Q, QN;
input D, SI, SE, CK, RN;
supply1 xSN;
supply1 dSN;

  udp_dff_PWR I0 (n0, n1, CK, RN, xSN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFRXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSHQX1 (Q, CK, D, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN;
supply1 xRN;
supply1 dRN;

  udp_dff_PWR I0 (n0, n1, CK, xRN, SN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFSHQX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSHQX2 (Q, CK, D, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN;
supply1 xRN;
supply1 dRN;

  udp_dff_PWR I0 (n0, n1, CK, xRN, SN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFSHQX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSHQX4 (Q, CK, D, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN;
supply1 xRN;
supply1 dRN;

  udp_dff_PWR I0 (n0, n1, CK, xRN, SN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFSHQX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSHQXL (Q, CK, D, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN;
supply1 xRN;
supply1 dRN;

  udp_dff_PWR I0 (n0, n1, CK, xRN, SN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFSHQXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRHQX1 (Q, CK, D, RN, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN, RN;
  udp_dff_PWR I0 (n0, n1, CK, RN, SN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFSRHQX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRHQX2 (Q, CK, D, RN, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN, RN;
  udp_dff_PWR I0 (n0, n1, CK, RN, SN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFSRHQX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRHQX4 (Q, CK, D, RN, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN, RN;
  udp_dff_PWR I0 (n0, n1, CK, RN, SN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFSRHQX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRHQXL (Q, CK, D, RN, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN, RN;
  udp_dff_PWR I0 (n0, n1, CK, RN, SN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
endmodule // SDFFSRHQXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRX1 (Q, QN, CK, D, RN, SE, SI, SN);
output Q, QN;
input D, SI, SE, CK, SN, RN;
  udp_dff_PWR I0 (n0, n1, CK, RN, SN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFSRX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRX2 (Q, QN, CK, D, RN, SE, SI, SN);
output Q, QN;
input D, SI, SE, CK, SN, RN;
  udp_dff_PWR I0 (n0, n1, CK, RN, SN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFSRX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRX4 (Q, QN, CK, D, RN, SE, SI, SN);
output Q, QN;
input D, SI, SE, CK, SN, RN;
  udp_dff_PWR I0 (n0, n1, CK, RN, SN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFSRX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRXL (Q, QN, CK, D, RN, SE, SI, SN);
output Q, QN;
input D, SI, SE, CK, SN, RN;
  udp_dff_PWR I0 (n0, n1, CK, RN, SN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFSRXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSX1 (Q, QN, CK, D, SE, SI, SN);
output Q, QN;
input D, SI, SE, CK, SN;
supply1 xRN;
supply1 dRN;

  udp_dff_PWR I0 (n0, n1, CK, xRN, SN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFSX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSX2 (Q, QN, CK, D, SE, SI, SN);
output Q, QN;
input D, SI, SE, CK, SN;
supply1 xRN;
supply1 dRN;

  udp_dff_PWR I0 (n0, n1, CK, xRN, SN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFSX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSX4 (Q, QN, CK, D, SE, SI, SN);
output Q, QN;
input D, SI, SE, CK, SN;
supply1 xRN;
supply1 dRN;

  udp_dff_PWR I0 (n0, n1, CK, xRN, SN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFSX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSXL (Q, QN, CK, D, SE, SI, SN);
output Q, QN;
input D, SI, SE, CK, SN;
supply1 xRN;
supply1 dRN;

  udp_dff_PWR I0 (n0, n1, CK, xRN, SN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFSXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFTRX1 (Q, QN, CK, D, RN, SE, SI);
output Q, QN;
input D, SI, SE, CK, RN;
supply1 xSN;
supply1 dSN;

   udp_sedfft_PWR I0 (n0, D, CK, RN, SI, SE, 1'b1, 1'b1, 1'b0, 1'b1);
   buf        `ARM_UD_SEQ I1 (Q, n0);
   not        `ARM_UD_SEQ I2 (QN, n0);
endmodule // SDFFTRX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFTRX2 (Q, QN, CK, D, RN, SE, SI);
output Q, QN;
input D, SI, SE, CK, RN;
supply1 xSN;
supply1 dSN;

   udp_sedfft_PWR I0 (n0, D, CK, RN, SI, SE, 1'b1, 1'b1, 1'b0, 1'b1);
   buf        `ARM_UD_SEQ I1 (Q, n0);
   not        `ARM_UD_SEQ I2 (QN, n0);
endmodule // SDFFTRX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFTRX4 (Q, QN, CK, D, RN, SE, SI);
output Q, QN;
input D, SI, SE, CK, RN;
supply1 xSN;
supply1 dSN;

   udp_sedfft_PWR I0 (n0, D, CK, RN, SI, SE, 1'b1, 1'b1, 1'b0, 1'b1);
   buf        `ARM_UD_SEQ I1 (Q, n0);
   not        `ARM_UD_SEQ I2 (QN, n0);
endmodule // SDFFTRX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFTRXL (Q, QN, CK, D, RN, SE, SI);
output Q, QN;
input D, SI, SE, CK, RN;
supply1 xSN;
supply1 dSN;

   udp_sedfft_PWR I0 (n0, D, CK, RN, SI, SE, 1'b1, 1'b1, 1'b0, 1'b1);
   buf        `ARM_UD_SEQ I1 (Q, n0);
   not        `ARM_UD_SEQ I2 (QN, n0);
endmodule // SDFFTRXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFX1 (Q, QN, CK, D, SE, SI);
output Q, QN;
input D, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  udp_dff_PWR I0 (n0, n1, CK, xRN, xSN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFX2 (Q, QN, CK, D, SE, SI);
output Q, QN;
input D, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  udp_dff_PWR I0 (n0, n1, CK, xRN, xSN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFX4 (Q, QN, CK, D, SE, SI);
output Q, QN;
input D, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  udp_dff_PWR I0 (n0, n1, CK, xRN, xSN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFXL (Q, QN, CK, D, SE, SI);
output Q, QN;
input D, SI, SE, CK;
supply1 xRN, xSN;
supply1 dRN, dSN;
  udp_dff_PWR I0 (n0, n1, CK, xRN, xSN, 1'b1, 1'b0, 1'b1);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     `ARM_UD_SEQ I2 (Q, n0);
  not     `ARM_UD_SEQ I72 (QN, n0);
endmodule // SDFFXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SEDFFHQX1 (Q, CK, D, E, SE, SI);
output Q;
input D, CK, E, SE, SI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR I0 (n0, D, CK, xRN, SI, SE, E, 1'b1, 1'b0, 1'b1);
   buf       `ARM_UD_SEQ I1 (Q, n0);
endmodule // SEDFFHQX1
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFHQX2 (Q, CK, D, E, SE, SI);
output Q;
input D, CK, E, SE, SI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR I0 (n0, D, CK, xRN, SI, SE, E, 1'b1, 1'b0, 1'b1);
   buf       `ARM_UD_SEQ I1 (Q, n0);
endmodule // SEDFFHQX2
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFHQX4 (Q, CK, D, E, SE, SI);
output Q;
input D, CK, E, SE, SI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR I0 (n0, D, CK, xRN, SI, SE, E, 1'b1, 1'b0, 1'b1);
   buf       `ARM_UD_SEQ I1 (Q, n0);
endmodule // SEDFFHQX4
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFHQXL (Q, CK, D, E, SE, SI);
output Q;
input D, CK, E, SE, SI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR I0 (n0, D, CK, xRN, SI, SE, E, 1'b1, 1'b0, 1'b1);
   buf       `ARM_UD_SEQ I1 (Q, n0);
endmodule // SEDFFHQXL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFTRX1 (Q, QN, CK, D, E, RN, SE, SI);
output Q, QN;
input D, CK, E, SE, SI, RN;
supply1 xSN;
supply1 dSN;

   udp_sedfft_PWR I0 (n0, D, CK, RN, SI, SE, E, 1'b1, 1'b0, 1'b1);
   buf        `ARM_UD_SEQ I1 (Q, n0);
   not        `ARM_UD_SEQ I2 (QN, n0);
endmodule // SEDFFTRX1
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFTRX2 (Q, QN, CK, D, E, RN, SE, SI);
output Q, QN;
input D, CK, E, SE, SI, RN;
supply1 xSN;
supply1 dSN;

   udp_sedfft_PWR I0 (n0, D, CK, RN, SI, SE, E, 1'b1, 1'b0, 1'b1);
   buf        `ARM_UD_SEQ I1 (Q, n0);
   not        `ARM_UD_SEQ I2 (QN, n0);
endmodule // SEDFFTRX2
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFTRX4 (Q, QN, CK, D, E, RN, SE, SI);
output Q, QN;
input D, CK, E, SE, SI, RN;
supply1 xSN;
supply1 dSN;

   udp_sedfft_PWR I0 (n0, D, CK, RN, SI, SE, E, 1'b1, 1'b0, 1'b1);
   buf        `ARM_UD_SEQ I1 (Q, n0);
   not        `ARM_UD_SEQ I2 (QN, n0);
endmodule // SEDFFTRX4
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFTRXL (Q, QN, CK, D, E, RN, SE, SI);
output Q, QN;
input D, CK, E, SE, SI, RN;
supply1 xSN;
supply1 dSN;

   udp_sedfft_PWR I0 (n0, D, CK, RN, SI, SE, E, 1'b1, 1'b0, 1'b1);
   buf        `ARM_UD_SEQ I1 (Q, n0);
   not        `ARM_UD_SEQ I2 (QN, n0);
endmodule // SEDFFTRXL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFX1 (Q, QN, CK, D, E, SE, SI);
output Q, QN;
input D, CK, E, SE, SI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR I0 (n0, D, CK, xRN, SI, SE, E, 1'b1, 1'b0, 1'b1); 
  buf     `ARM_UD_SEQ I1 (Q, n0);  
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // SEDFFX1
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFX2 (Q, QN, CK, D, E, SE, SI);
output Q, QN;
input D, CK, E, SE, SI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR I0 (n0, D, CK, xRN, SI, SE, E, 1'b1, 1'b0, 1'b1); 
  buf     `ARM_UD_SEQ I1 (Q, n0);  
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // SEDFFX2
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFX4 (Q, QN, CK, D, E, SE, SI);
output Q, QN;
input D, CK, E, SE, SI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR I0 (n0, D, CK, xRN, SI, SE, E, 1'b1, 1'b0, 1'b1); 
  buf     `ARM_UD_SEQ I1 (Q, n0);  
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // SEDFFX4
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFXL (Q, QN, CK, D, E, SE, SI);
output Q, QN;
input D, CK, E, SE, SI;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR I0 (n0, D, CK, xRN, SI, SE, E, 1'b1, 1'b0, 1'b1); 
  buf     `ARM_UD_SEQ I1 (Q, n0);  
  not     `ARM_UD_SEQ I2 (QN, n0);
endmodule // SEDFFXL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module TBUFIX1 (Y, A, OE);
output Y;
input A, OE;

  notif1 `ARM_UD_DP I0(Y, A, OE);

endmodule // TBUFIX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFIX12 (Y, A, OE);
output Y;
input A, OE;

  notif1 `ARM_UD_DP I0(Y, A, OE);

endmodule // TBUFIX12
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFIX16 (Y, A, OE);
output Y;
input A, OE;

  notif1 `ARM_UD_DP I0(Y, A, OE);

endmodule // TBUFIX16
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFIX2 (Y, A, OE);
output Y;
input A, OE;

  notif1 `ARM_UD_DP I0(Y, A, OE);

endmodule // TBUFIX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFIX20 (Y, A, OE);
output Y;
input A, OE;

  notif1 `ARM_UD_DP I0(Y, A, OE);

endmodule // TBUFIX20
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFIX3 (Y, A, OE);
output Y;
input A, OE;

  notif1 `ARM_UD_DP I0(Y, A, OE);

endmodule // TBUFIX3
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFIX4 (Y, A, OE);
output Y;
input A, OE;

  notif1 `ARM_UD_DP I0(Y, A, OE);

endmodule // TBUFIX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFIX8 (Y, A, OE);
output Y;
input A, OE;

  notif1 `ARM_UD_DP I0(Y, A, OE);

endmodule // TBUFIX8
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFIXL (Y, A, OE);
output Y;
input A, OE;

  notif1 `ARM_UD_DP I0(Y, A, OE);

endmodule // TBUFIXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFX1 (Y, A, OE);
output Y;
input A, OE;

  bufif1 `ARM_UD_DP I0(Y, A, OE);

endmodule // TBUFX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFX12 (Y, A, OE);
output Y;
input A, OE;

  bufif1 `ARM_UD_DP I0(Y, A, OE);

endmodule // TBUFX12
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFX16 (Y, A, OE);
output Y;
input A, OE;

  bufif1 `ARM_UD_DP I0(Y, A, OE);

endmodule // TBUFX16
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFX2 (Y, A, OE);
output Y;
input A, OE;

  bufif1 `ARM_UD_DP I0(Y, A, OE);

endmodule // TBUFX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFX20 (Y, A, OE);
output Y;
input A, OE;

  bufif1 `ARM_UD_DP I0(Y, A, OE);

endmodule // TBUFX20
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFX3 (Y, A, OE);
output Y;
input A, OE;

  bufif1 `ARM_UD_DP I0(Y, A, OE);

endmodule // TBUFX3
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFX4 (Y, A, OE);
output Y;
input A, OE;

  bufif1 `ARM_UD_DP I0(Y, A, OE);

endmodule // TBUFX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFX8 (Y, A, OE);
output Y;
input A, OE;

  bufif1 `ARM_UD_DP I0(Y, A, OE);

endmodule // TBUFX8
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFXL (Y, A, OE);
output Y;
input A, OE;

  bufif1 `ARM_UD_DP I0(Y, A, OE);

endmodule // TBUFXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TIEHI (Y);
output Y;

  buf I0(Y, 1'b1);

endmodule // TIEHI
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TIELO (Y);
output Y;

  buf I0(Y, 1'b0);

endmodule // TIELO
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATCOX1 (ECKN, CKN, E);
output ECKN;
input  E, CKN;

supply1 R, S;

  not      I0 (nclk,CKN);
  udp_tlat_PWR I1 (n0, E, nclk, R, S, 1'b1, 1'b0, 1'b1);
  not      I2 (nn0,n0);
  or       `ARM_UD_CP I3 (ECKN, nn0, CKN);

endmodule // TLATCOX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATCOX2 (ECKN, CKN, E);
output ECKN;
input  E, CKN;

supply1 R, S;

  not      I0 (nclk,CKN);
  udp_tlat_PWR I1 (n0, E, nclk, R, S, 1'b1, 1'b0, 1'b1);
  not      I2 (nn0,n0);
  or       `ARM_UD_CP I3 (ECKN, nn0, CKN);

endmodule // TLATCOX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATCOX3 (ECKN, CKN, E);
output ECKN;
input  E, CKN;

supply1 R, S;

  not      I0 (nclk,CKN);
  udp_tlat_PWR I1 (n0, E, nclk, R, S, 1'b1, 1'b0, 1'b1);
  not      I2 (nn0,n0);
  or       `ARM_UD_CP I3 (ECKN, nn0, CKN);

endmodule // TLATCOX3
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATCOX4 (ECKN, CKN, E);
output ECKN;
input  E, CKN;

supply1 R, S;

  not      I0 (nclk,CKN);
  udp_tlat_PWR I1 (n0, E, nclk, R, S, 1'b1, 1'b0, 1'b1);
  not      I2 (nn0,n0);
  or       `ARM_UD_CP I3 (ECKN, nn0, CKN);

endmodule // TLATCOX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNCAX1 (ECK, CK, E);
output ECK;
input  E, CK;

supply1 R, S;

  udp_tlat_PWR I0 (n0, E, CK, R, S, 1'b1, 1'b0, 1'b1);
  and      `ARM_UD_CP I1 (ECK, n0, CK);

endmodule // TLATNCAX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNCAX2 (ECK, CK, E);
output ECK;
input  E, CK;

supply1 R, S;

  udp_tlat_PWR I0 (n0, E, CK, R, S, 1'b1, 1'b0, 1'b1);
  and      `ARM_UD_CP I1 (ECK, n0, CK);

endmodule // TLATNCAX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNCAX3 (ECK, CK, E);
output ECK;
input  E, CK;

supply1 R, S;

  udp_tlat_PWR I0 (n0, E, CK, R, S, 1'b1, 1'b0, 1'b1);
  and      `ARM_UD_CP I1 (ECK, n0, CK);

endmodule // TLATNCAX3
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNCAX4 (ECK, CK, E);
output ECK;
input  E, CK;

supply1 R, S;

  udp_tlat_PWR I0 (n0, E, CK, R, S, 1'b1, 1'b0, 1'b1);
  and      `ARM_UD_CP I1 (ECK, n0, CK);

endmodule // TLATNCAX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNCAX6 (ECK, CK, E);
output ECK;
input  E, CK;

supply1 R, S;

  udp_tlat_PWR I0 (n0, E, CK, R, S, 1'b1, 1'b0, 1'b1);
  and      `ARM_UD_CP I1 (ECK, n0, CK);

endmodule // TLATNCAX6
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNCAX8 (ECK, CK, E);
output ECK;
input  E, CK;

supply1 R, S;

  udp_tlat_PWR I0 (n0, E, CK, R, S, 1'b1, 1'b0, 1'b1);
  and      `ARM_UD_CP I1 (ECK, n0, CK);

endmodule // TLATNCAX8
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNRX1 (Q, QN, D, GN, RN);
output  Q, QN;
input  D, GN, RN;
supply1 xSN;
supply1 dSN;


udp_tlat_PWR I0 (n0, D, GN, RN, xSN, 1'b1, 1'b0, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not      `ARM_UD_SEQ I2 (QN, n0);
endmodule // TLATNRX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNRX2 (Q, QN, D, GN, RN);
output  Q, QN;
input  D, GN, RN;
supply1 xSN;
supply1 dSN;


udp_tlat_PWR I0 (n0, D, GN, RN, xSN, 1'b1, 1'b0, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not      `ARM_UD_SEQ I2 (QN, n0);
endmodule // TLATNRX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNRX4 (Q, QN, D, GN, RN);
output  Q, QN;
input  D, GN, RN;
supply1 xSN;
supply1 dSN;


udp_tlat_PWR I0 (n0, D, GN, RN, xSN, 1'b1, 1'b0, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not      `ARM_UD_SEQ I2 (QN, n0);
endmodule // TLATNRX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNRXL (Q, QN, D, GN, RN);
output  Q, QN;
input  D, GN, RN;
supply1 xSN;
supply1 dSN;


udp_tlat_PWR I0 (n0, D, GN, RN, xSN, 1'b1, 1'b0, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not      `ARM_UD_SEQ I2 (QN, n0);
endmodule // TLATNRXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNSRX1 (Q, QN, D, GN, RN, SN);
output  Q, QN;
input  D, GN, RN, SN;


udp_tlat_PWR I0 (n0, D, GN, RN, SN, 1'b1, 1'b0, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not      `ARM_UD_SEQ I2 (QN, n0);
buf      I3 (clk, GN);
endmodule // TLATNSRX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNSRX2 (Q, QN, D, GN, RN, SN);
output  Q, QN;
input  D, GN, RN, SN;


udp_tlat_PWR I0 (n0, D, GN, RN, SN, 1'b1, 1'b0, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not      `ARM_UD_SEQ I2 (QN, n0);
buf      I3 (clk, GN);
endmodule // TLATNSRX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNSRX4 (Q, QN, D, GN, RN, SN);
output  Q, QN;
input  D, GN, RN, SN;


udp_tlat_PWR I0 (n0, D, GN, RN, SN, 1'b1, 1'b0, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not      `ARM_UD_SEQ I2 (QN, n0);
buf      I3 (clk, GN);
endmodule // TLATNSRX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNSRXL (Q, QN, D, GN, RN, SN);
output  Q, QN;
input  D, GN, RN, SN;


udp_tlat_PWR I0 (n0, D, GN, RN, SN, 1'b1, 1'b0, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not      `ARM_UD_SEQ I2 (QN, n0);
buf      I3 (clk, GN);
endmodule // TLATNSRXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNSX1 (Q, QN, D, GN, SN);
output  Q, QN;
input  D, GN, SN;
supply1 xRN;
supply1 dRN;


udp_tlat_PWR I0 (n0, D, GN, xRN, SN, 1'b1, 1'b0, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not      `ARM_UD_SEQ I2 (QN, n0);
endmodule // TLATNSX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNSX2 (Q, QN, D, GN, SN);
output  Q, QN;
input  D, GN, SN;
supply1 xRN;
supply1 dRN;


udp_tlat_PWR I0 (n0, D, GN, xRN, SN, 1'b1, 1'b0, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not      `ARM_UD_SEQ I2 (QN, n0);
endmodule // TLATNSX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNSX4 (Q, QN, D, GN, SN);
output  Q, QN;
input  D, GN, SN;
supply1 xRN;
supply1 dRN;


udp_tlat_PWR I0 (n0, D, GN, xRN, SN, 1'b1, 1'b0, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not      `ARM_UD_SEQ I2 (QN, n0);
endmodule // TLATNSX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNSXL (Q, QN, D, GN, SN);
output  Q, QN;
input  D, GN, SN;
supply1 xRN;
supply1 dRN;


udp_tlat_PWR I0 (n0, D, GN, xRN, SN, 1'b1, 1'b0, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not      `ARM_UD_SEQ I2 (QN, n0);
endmodule // TLATNSXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNTSCAX1 (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR I1 (n0, n1, CK, R, S, 1'b1, 1'b0, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // TLATNTSCAX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNTSCAX2 (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR I1 (n0, n1, CK, R, S, 1'b1, 1'b0, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // TLATNTSCAX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNTSCAX3 (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR I1 (n0, n1, CK, R, S, 1'b1, 1'b0, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // TLATNTSCAX3
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNTSCAX4 (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR I1 (n0, n1, CK, R, S, 1'b1, 1'b0, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // TLATNTSCAX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNTSCAX6 (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR I1 (n0, n1, CK, R, S, 1'b1, 1'b0, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // TLATNTSCAX6
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNTSCAX8 (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR I1 (n0, n1, CK, R, S, 1'b1, 1'b0, 1'b1);
  and      `ARM_UD_CP I2 (ECK, n0, CK);

endmodule // TLATNTSCAX8
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNX1 (Q, QN, D, GN);
output  Q, QN;
input  D, GN;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR I0 (n0, D, GN, xRN, xSN, 1'b1, 1'b0, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not      `ARM_UD_SEQ I2 (QN, n0);
buf      I3 (clk, GN);
endmodule // TLATNX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNX2 (Q, QN, D, GN);
output  Q, QN;
input  D, GN;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR I0 (n0, D, GN, xRN, xSN, 1'b1, 1'b0, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not      `ARM_UD_SEQ I2 (QN, n0);
buf      I3 (clk, GN);
endmodule // TLATNX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNX4 (Q, QN, D, GN);
output  Q, QN;
input  D, GN;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR I0 (n0, D, GN, xRN, xSN, 1'b1, 1'b0, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not      `ARM_UD_SEQ I2 (QN, n0);
buf      I3 (clk, GN);
endmodule // TLATNX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNXL (Q, QN, D, GN);
output  Q, QN;
input  D, GN;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR I0 (n0, D, GN, xRN, xSN, 1'b1, 1'b0, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not      `ARM_UD_SEQ I2 (QN, n0);
buf      I3 (clk, GN);
endmodule // TLATNXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATRX1 (Q, QN, D, G, RN);
output  Q, QN;
input  D, G, RN;
supply1 xSN;
supply1 dSN;


udp_tlat_PWR I0 (n0, D, clk, RN, xSN, 1'b1, 1'b0, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not      `ARM_UD_SEQ I2 (QN, n0);
not  I3(clk,G);
endmodule // TLATRX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATRX2 (Q, QN, D, G, RN);
output  Q, QN;
input  D, G, RN;
supply1 xSN;
supply1 dSN;


udp_tlat_PWR I0 (n0, D, clk, RN, xSN, 1'b1, 1'b0, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not      `ARM_UD_SEQ I2 (QN, n0);
not  I3(clk,G);
endmodule // TLATRX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATRX4 (Q, QN, D, G, RN);
output  Q, QN;
input  D, G, RN;
supply1 xSN;
supply1 dSN;


udp_tlat_PWR I0 (n0, D, clk, RN, xSN, 1'b1, 1'b0, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not      `ARM_UD_SEQ I2 (QN, n0);
not  I3(clk,G);
endmodule // TLATRX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATRXL (Q, QN, D, G, RN);
output  Q, QN;
input  D, G, RN;
supply1 xSN;
supply1 dSN;


udp_tlat_PWR I0 (n0, D, clk, RN, xSN, 1'b1, 1'b0, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not      `ARM_UD_SEQ I2 (QN, n0);
not  I3(clk,G);
endmodule // TLATRXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATSRX1 (Q, QN, D, G, RN, SN);
output  Q, QN;
input  D, G, SN, RN;


udp_tlat_PWR I0 (n0, D, clk, RN, SN, 1'b1, 1'b0, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not      `ARM_UD_SEQ I2 (QN, n0);
not  I3(clk,G);
endmodule // TLATSRX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATSRX2 (Q, QN, D, G, RN, SN);
output  Q, QN;
input  D, G, SN, RN;


udp_tlat_PWR I0 (n0, D, clk, RN, SN, 1'b1, 1'b0, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not      `ARM_UD_SEQ I2 (QN, n0);
not  I3(clk,G);
endmodule // TLATSRX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATSRX4 (Q, QN, D, G, RN, SN);
output  Q, QN;
input  D, G, SN, RN;


udp_tlat_PWR I0 (n0, D, clk, RN, SN, 1'b1, 1'b0, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not      `ARM_UD_SEQ I2 (QN, n0);
not  I3(clk,G);
endmodule // TLATSRX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATSRXL (Q, QN, D, G, RN, SN);
output  Q, QN;
input  D, G, SN, RN;


udp_tlat_PWR I0 (n0, D, clk, RN, SN, 1'b1, 1'b0, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not      `ARM_UD_SEQ I2 (QN, n0);
not  I3(clk,G);
endmodule // TLATSRXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATSX1 (Q, QN, D, G, SN);
output  Q, QN;
input  D, G, SN;
supply1 xRN;
supply1 dRN;


udp_tlat_PWR I0 (n0, D, clk, xRN, SN, 1'b1, 1'b0, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not      `ARM_UD_SEQ I2 (QN, n0);
not  I3(clk,G);
endmodule // TLATSX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATSX2 (Q, QN, D, G, SN);
output  Q, QN;
input  D, G, SN;
supply1 xRN;
supply1 dRN;


udp_tlat_PWR I0 (n0, D, clk, xRN, SN, 1'b1, 1'b0, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not      `ARM_UD_SEQ I2 (QN, n0);
not  I3(clk,G);
endmodule // TLATSX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATSX4 (Q, QN, D, G, SN);
output  Q, QN;
input  D, G, SN;
supply1 xRN;
supply1 dRN;


udp_tlat_PWR I0 (n0, D, clk, xRN, SN, 1'b1, 1'b0, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not      `ARM_UD_SEQ I2 (QN, n0);
not  I3(clk,G);
endmodule // TLATSX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATSXL (Q, QN, D, G, SN);
output  Q, QN;
input  D, G, SN;
supply1 xRN;
supply1 dRN;


udp_tlat_PWR I0 (n0, D, clk, xRN, SN, 1'b1, 1'b0, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not      `ARM_UD_SEQ I2 (QN, n0);
not  I3(clk,G);
endmodule // TLATSXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATTSCOX1 (ECKN, CKN, E, SE);
output ECKN;
input  E, SE, CKN;

supply1 R, S;

  not      I0 (nclk,CKN);
  or       I1 (n1, SE, E);
  udp_tlat_PWR I2 (n0, n1, nclk, R, S, 1'b1, 1'b0, 1'b1);
  not      I3 (nn0,n0);
  or       `ARM_UD_CP I4 (ECKN, nn0, CKN);

endmodule // TLATTSCOX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATTSCOX2 (ECKN, CKN, E, SE);
output ECKN;
input  E, SE, CKN;

supply1 R, S;

  not      I0 (nclk,CKN);
  or       I1 (n1, SE, E);
  udp_tlat_PWR I2 (n0, n1, nclk, R, S, 1'b1, 1'b0, 1'b1);
  not      I3 (nn0,n0);
  or       `ARM_UD_CP I4 (ECKN, nn0, CKN);

endmodule // TLATTSCOX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATTSCOX3 (ECKN, CKN, E, SE);
output ECKN;
input  E, SE, CKN;

supply1 R, S;

  not      I0 (nclk,CKN);
  or       I1 (n1, SE, E);
  udp_tlat_PWR I2 (n0, n1, nclk, R, S, 1'b1, 1'b0, 1'b1);
  not      I3 (nn0,n0);
  or       `ARM_UD_CP I4 (ECKN, nn0, CKN);

endmodule // TLATTSCOX3
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATTSCOX4 (ECKN, CKN, E, SE);
output ECKN;
input  E, SE, CKN;

supply1 R, S;

  not      I0 (nclk,CKN);
  or       I1 (n1, SE, E);
  udp_tlat_PWR I2 (n0, n1, nclk, R, S, 1'b1, 1'b0, 1'b1);
  not      I3 (nn0,n0);
  or       `ARM_UD_CP I4 (ECKN, nn0, CKN);

endmodule // TLATTSCOX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATX1 (Q, QN, D, G);
output  Q, QN;
input  D, G;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not      `ARM_UD_SEQ I2 (QN, n0);
not  I3(clk,G);
endmodule // TLATX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATX2 (Q, QN, D, G);
output  Q, QN;
input  D, G;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not      `ARM_UD_SEQ I2 (QN, n0);
not  I3(clk,G);
endmodule // TLATX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATX4 (Q, QN, D, G);
output  Q, QN;
input  D, G;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not      `ARM_UD_SEQ I2 (QN, n0);
not  I3(clk,G);
endmodule // TLATX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATXL (Q, QN, D, G);
output  Q, QN;
input  D, G;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, 1'b1);
buf      `ARM_UD_SEQ I1 (Q, n0);
not      `ARM_UD_SEQ I2 (QN, n0);
not  I3(clk,G);
endmodule // TLATXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TTLATX1 (Q, D, G, OE);
output Q;
input  D, G, OE;
supply1 RN, SN;
supply1 xRN, xSN;
supply1 dRN, dSN;

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, 1'b1);
bufif1   `ARM_UD_SEQ I1 (Q, n0, OE);
not  I3(clk,G);
endmodule // TTLATX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TTLATX2 (Q, D, G, OE);
output Q;
input  D, G, OE;
supply1 RN, SN;
supply1 xRN, xSN;
supply1 dRN, dSN;

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, 1'b1);
bufif1   `ARM_UD_SEQ I1 (Q, n0, OE);
not  I3(clk,G);
endmodule // TTLATX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TTLATX4 (Q, D, G, OE);
output Q;
input  D, G, OE;
supply1 RN, SN;
supply1 xRN, xSN;
supply1 dRN, dSN;

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, 1'b1);
bufif1   `ARM_UD_SEQ I1 (Q, n0, OE);
not  I3(clk,G);
endmodule // TTLATX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TTLATXL (Q, D, G, OE);
output Q;
input  D, G, OE;
supply1 RN, SN;
supply1 xRN, xSN;
supply1 dRN, dSN;

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, 1'b1);
bufif1   `ARM_UD_SEQ I1 (Q, n0, OE);
not  I3(clk,G);
endmodule // TTLATXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2X1 (Y, A, B);
output Y;
input A, B;

  xnor `ARM_UD_DP I0(Y, A, B);

endmodule // XNOR2X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2X2 (Y, A, B);
output Y;
input A, B;

  xnor `ARM_UD_DP I0(Y, A, B);

endmodule // XNOR2X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2X4 (Y, A, B);
output Y;
input A, B;

  xnor `ARM_UD_DP I0(Y, A, B);

endmodule // XNOR2X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2XL (Y, A, B);
output Y;
input A, B;

  xnor `ARM_UD_DP I0(Y, A, B);

endmodule // XNOR2XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3X2 (Y, A, B, C);
output Y;
input A, B, C;

  xnor `ARM_UD_DP I0(Y, A, B, C);

endmodule // XNOR3X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3X4 (Y, A, B, C);
output Y;
input A, B, C;

  xnor `ARM_UD_DP I0(Y, A, B, C);

endmodule // XNOR3X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2X1 (Y, A, B);
output Y;
input A, B;

  xor `ARM_UD_DP I0(Y, A, B);

endmodule // XOR2X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2X2 (Y, A, B);
output Y;
input A, B;

  xor `ARM_UD_DP I0(Y, A, B);

endmodule // XOR2X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2X4 (Y, A, B);
output Y;
input A, B;

  xor `ARM_UD_DP I0(Y, A, B);

endmodule // XOR2X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2XL (Y, A, B);
output Y;
input A, B;

  xor `ARM_UD_DP I0(Y, A, B);

endmodule // XOR2XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3X2 (Y, A, B, C);
output Y;
input A, B, C;

  xor `ARM_UD_DP I0(Y, A, B, C);

endmodule // XOR3X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3X4 (Y, A, B, C);
output Y;
input A, B, C;

  xor `ARM_UD_DP I0(Y, A, B, C);

endmodule // XOR3X4
`endcelldefine
`else

`timescale 1ns/1ps
`define ARM_PROP_DELAY 		1.0
`define ARM_INVALID_DELAY 	1.0

`define ARM_PERIOD 			1.0
`define ARM_WIDTH 			1.0
`define ARM_SETUP_TIME 		1.0
`define ARM_HOLD_TIME 		0.5
`define ARM_RECOVERY_TIME 	1.0
`define ARM_REMOVAL_TIME 	0.5
`define ARM_WIDTH_THD 		0.0

`ifdef POWER_PINS
`timescale 1ns/1ps
`celldefine
module ADDFHX1 (CO, S, VDD, VSS, A, B, CI);
inout VDD, VSS;
output S, CO;
input A, B, CI;
  xor I0(S_temp, A, B, CI);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? S_temp : 1'bx;
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(cout_temp, a_and_b, a_and_ci, b_and_ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFHX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFHX2 (CO, S, VDD, VSS, A, B, CI);
inout VDD, VSS;
output S, CO;
input A, B, CI;
  xor I0(S_temp, A, B, CI);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? S_temp : 1'bx;
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(cout_temp, a_and_b, a_and_ci, b_and_ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFHX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFHX4 (CO, S, VDD, VSS, A, B, CI);
inout VDD, VSS;
output S, CO;
input A, B, CI;
  xor I0(S_temp, A, B, CI);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? S_temp : 1'bx;
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(cout_temp, a_and_b, a_and_ci, b_and_ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFHX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFHXL (CO, S, VDD, VSS, A, B, CI);
inout VDD, VSS;
output S, CO;
input A, B, CI;
  xor I0(S_temp, A, B, CI);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? S_temp : 1'bx;
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(cout_temp, a_and_b, a_and_ci, b_and_ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFHXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFX1 (CO, S, VDD, VSS, A, B, CI);
inout VDD, VSS;
output S, CO;
input A, B, CI;
  xor I0(sum_temp, A, B, CI);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(cout_temp, a_and_b, a_and_ci, b_and_ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFX2 (CO, S, VDD, VSS, A, B, CI);
inout VDD, VSS;
output S, CO;
input A, B, CI;
  xor I0(sum_temp, A, B, CI);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(cout_temp, a_and_b, a_and_ci, b_and_ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFX4 (CO, S, VDD, VSS, A, B, CI);
inout VDD, VSS;
output S, CO;
input A, B, CI;
  xor I0(sum_temp, A, B, CI);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(cout_temp, a_and_b, a_and_ci, b_and_ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFXL (CO, S, VDD, VSS, A, B, CI);
inout VDD, VSS;
output S, CO;
input A, B, CI;
  xor I0(sum_temp, A, B, CI);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(cout_temp, a_and_b, a_and_ci, b_and_ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDHX1 (CO, S, VDD, VSS, A, B);
inout VDD, VSS;
output S, CO;
input A, B;
  xor I0(sum_temp, A, B);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I1(cout_temp, A, B);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDHX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDHX2 (CO, S, VDD, VSS, A, B);
inout VDD, VSS;
output S, CO;
input A, B;
  xor I0(sum_temp, A, B);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I1(cout_temp, A, B);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDHX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDHX4 (CO, S, VDD, VSS, A, B);
inout VDD, VSS;
output S, CO;
input A, B;
  xor I0(sum_temp, A, B);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I1(cout_temp, A, B);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDHX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDHXL (CO, S, VDD, VSS, A, B);
inout VDD, VSS;
output S, CO;
input A, B;
  xor I0(sum_temp, A, B);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I1(cout_temp, A, B);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDHXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AFCSHCINX2 (CO0, CO1, S, VDD, VSS, A, B, CI0N, CI1N, CS);
inout VDD, VSS;
output S, CO0, CO1;
input A, B, CI0N, CI1N, CS;
  not I0 (cin1, CI1N);
  not I1 (cin0, CI0N);
  xor I2 (s1, A, B, cin1);
  xor I3 (s2, A, B, cin0);
  and I4 (s3, CS, s1);
  not I5 (csn, CS);
  and I6 (s4, csn, s2);
  or I7 (sum_temp, s3, s4);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I8 (a_and_b, A, B);
  and I9 (a_and_ci0, A, cin0);
  and I10 (b_and_ci0, B, cin0);
  or I11 (cout0_temp, a_and_b, a_and_ci0, b_and_ci0);
  assign CO0 = ((VDD === 1'b1) && (VSS === 1'b0))? cout0_temp : 1'bx;
  and I12 (a_and_ci1, A, cin1);
  and I13 (b_and_ci1, B, cin1);
  or I14 (cout1_temp, a_and_b, a_and_ci1, b_and_ci1);
  assign CO1 = ((VDD === 1'b1) && (VSS === 1'b0))? cout1_temp : 1'bx;


specify
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b0)
(A => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b1)
(A => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b0)
(A => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b1)
(A => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b0)
(A => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b1)
(A => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b0)
(A => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b1)
(A => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b0)
(B => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b1)
(B => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b0)
(B => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b1)
(B => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b0)
(B => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b1)
(B => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b0)
(B => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b1)
(B => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1N==1'b0 && CS==1'b0)
(CI0N => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1N==1'b0 && CS==1'b1)
(CI0N => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1N==1'b1 && CS==1'b0)
(CI0N => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1N==1'b1 && CS==1'b1)
(CI0N => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1N==1'b0 && CS==1'b0)
(CI0N => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1N==1'b0 && CS==1'b1)
(CI0N => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1N==1'b1 && CS==1'b0)
(CI0N => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1N==1'b1 && CS==1'b1)
(CI0N => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b0)
(A => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b1)
(A => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b0)
(A => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b1)
(A => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b0)
(A => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b1)
(A => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b0)
(A => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b1)
(A => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b0)
(B => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b1)
(B => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b0)
(B => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b1)
(B => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b0)
(B => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b1)
(B => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b0)
(B => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b1)
(B => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0N==1'b0 && CS==1'b0)
(CI1N => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0N==1'b0 && CS==1'b1)
(CI1N => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0N==1'b1 && CS==1'b0)
(CI1N => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0N==1'b1 && CS==1'b1)
(CI1N => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0N==1'b0 && CS==1'b0)
(CI1N => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0N==1'b0 && CS==1'b1)
(CI1N => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0N==1'b1 && CS==1'b0)
(CI1N => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0N==1'b1 && CS==1'b1)
(CI1N => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI1N==1'b0)
(CI0N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI1N==1'b1)
(CI0N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI1N==1'b0)
(CI0N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI1N==1'b1)
(CI0N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1N==1'b0)
(CI0N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1N==1'b1)
(CI0N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1N==1'b0)
(CI0N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1N==1'b1)
(CI0N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI0N==1'b0)
(CI1N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI0N==1'b1)
(CI1N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI0N==1'b0)
(CI1N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI0N==1'b1)
(CI1N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0N==1'b0)
(CI1N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0N==1'b1)
(CI1N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0N==1'b0)
(CI1N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0N==1'b1)
(CI1N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI0N==1'b0 && CI1N==1'b1)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0N==1'b1 && CI1N==1'b0)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0N==1'b1 && CI1N==1'b0)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI0N==1'b0 && CI1N==1'b1)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI0N==1'b1 && CI1N==1'b0)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0N==1'b0 && CI1N==1'b1)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0N==1'b0 && CI1N==1'b1)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI0N==1'b1 && CI1N==1'b0)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AFCSHCINX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AFCSHCINX4 (CO0, CO1, S, VDD, VSS, A, B, CI0N, CI1N, CS);
inout VDD, VSS;
output S, CO0, CO1;
input A, B, CI0N, CI1N, CS;
  not I0 (cin1, CI1N);
  not I1 (cin0, CI0N);
  xor I2 (s1, A, B, cin1);
  xor I3 (s2, A, B, cin0);
  and I4 (s3, CS, s1);
  not I5 (csn, CS);
  and I6 (s4, csn, s2);
  or I7 (sum_temp, s3, s4);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I8 (a_and_b, A, B);
  and I9 (a_and_ci0, A, cin0);
  and I10 (b_and_ci0, B, cin0);
  or I11 (cout0_temp, a_and_b, a_and_ci0, b_and_ci0);
  assign CO0 = ((VDD === 1'b1) && (VSS === 1'b0))? cout0_temp : 1'bx;
  and I12 (a_and_ci1, A, cin1);
  and I13 (b_and_ci1, B, cin1);
  or I14 (cout1_temp, a_and_b, a_and_ci1, b_and_ci1);
  assign CO1 = ((VDD === 1'b1) && (VSS === 1'b0))? cout1_temp : 1'bx;


specify
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b0)
(A => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b1)
(A => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b0)
(A => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b1)
(A => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b0)
(A => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b1)
(A => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b0)
(A => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b1)
(A => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b0)
(B => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b1)
(B => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b0)
(B => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b1)
(B => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b0)
(B => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b1)
(B => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b0)
(B => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b1)
(B => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1N==1'b0 && CS==1'b0)
(CI0N => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1N==1'b0 && CS==1'b1)
(CI0N => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1N==1'b1 && CS==1'b0)
(CI0N => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1N==1'b1 && CS==1'b1)
(CI0N => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1N==1'b0 && CS==1'b0)
(CI0N => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1N==1'b0 && CS==1'b1)
(CI0N => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1N==1'b1 && CS==1'b0)
(CI0N => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1N==1'b1 && CS==1'b1)
(CI0N => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b0)
(A => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b1)
(A => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b0)
(A => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b1)
(A => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b0)
(A => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b1)
(A => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b0)
(A => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b1)
(A => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b0)
(B => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b1)
(B => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b0)
(B => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b1)
(B => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b0)
(B => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b1)
(B => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b0)
(B => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b1)
(B => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0N==1'b0 && CS==1'b0)
(CI1N => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0N==1'b0 && CS==1'b1)
(CI1N => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0N==1'b1 && CS==1'b0)
(CI1N => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0N==1'b1 && CS==1'b1)
(CI1N => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0N==1'b0 && CS==1'b0)
(CI1N => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0N==1'b0 && CS==1'b1)
(CI1N => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0N==1'b1 && CS==1'b0)
(CI1N => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0N==1'b1 && CS==1'b1)
(CI1N => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI1N==1'b0)
(CI0N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI1N==1'b1)
(CI0N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI1N==1'b0)
(CI0N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI1N==1'b1)
(CI0N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1N==1'b0)
(CI0N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1N==1'b1)
(CI0N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1N==1'b0)
(CI0N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1N==1'b1)
(CI0N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI0N==1'b0)
(CI1N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI0N==1'b1)
(CI1N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI0N==1'b0)
(CI1N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI0N==1'b1)
(CI1N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0N==1'b0)
(CI1N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0N==1'b1)
(CI1N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0N==1'b0)
(CI1N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0N==1'b1)
(CI1N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI0N==1'b0 && CI1N==1'b1)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0N==1'b1 && CI1N==1'b0)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0N==1'b1 && CI1N==1'b0)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI0N==1'b0 && CI1N==1'b1)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI0N==1'b1 && CI1N==1'b0)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0N==1'b0 && CI1N==1'b1)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0N==1'b0 && CI1N==1'b1)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI0N==1'b1 && CI1N==1'b0)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AFCSHCINX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AFCSHCONX2 (CO0N, CO1N, S, VDD, VSS, A, B, CI0, CI1, CS);
inout VDD, VSS;
output S, CO0N, CO1N;
input A, B, CI0, CI1, CS;
  xor I2 (s1, A, B, CI1);
  xor I3 (s2, A, B, CI0);
  and I4 (s3, CS, s1);
  not I5 (csn, CS);
  and I6 (s4, csn, s2);
  or I7 (sum_temp, s3, s4);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I8 (a_and_b, A, B);
  and I9 (a_and_ci0, A, CI0);
  and I10 (b_and_ci0, B, CI0);
  or I11 (cout0, a_and_b, a_and_ci0, b_and_ci0);
  and I12 (a_and_ci1, A, CI1);
  and I13 (b_and_ci1, B, CI1);
  or I14 (cout1, a_and_b, a_and_ci1, b_and_ci1);
  not I15 (cout0n_temp, cout0);
  assign CO0N = ((VDD === 1'b1) && (VSS === 1'b0))? cout0n_temp : 1'bx;
  not I16 (cout1n_temp, cout1);
  assign CO1N = ((VDD === 1'b1) && (VSS === 1'b0))? cout1n_temp : 1'bx;


specify
if (B==1'b0 && CI0==1'b1 && CI1==1'b0 && CS==1'b0)
(A => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b0 && CS==1'b1)
(A => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b0)
(A => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b1)
(A => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b0)
(A => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b1)
(A => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b1 && CS==1'b0)
(A => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b1 && CS==1'b1)
(A => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b0 && CS==1'b0)
(B => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b0 && CS==1'b1)
(B => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b0)
(B => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b1)
(B => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b0)
(B => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b1)
(B => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b1 && CS==1'b0)
(B => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b1 && CS==1'b1)
(B => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1==1'b0 && CS==1'b0)
(CI0 => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1==1'b0 && CS==1'b1)
(CI0 => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1==1'b1 && CS==1'b0)
(CI0 => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1==1'b1 && CS==1'b1)
(CI0 => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1==1'b0 && CS==1'b0)
(CI0 => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1==1'b0 && CS==1'b1)
(CI0 => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1==1'b1 && CS==1'b0)
(CI0 => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1==1'b1 && CS==1'b1)
(CI0 => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b0 && CI1==1'b1 && CS==1'b0)
(A => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b0 && CI1==1'b1 && CS==1'b1)
(A => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b0)
(A => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b1)
(A => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b0)
(A => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b1)
(A => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b1 && CI1==1'b0 && CS==1'b0)
(A => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b1 && CI1==1'b0 && CS==1'b1)
(A => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b0 && CI1==1'b1 && CS==1'b0)
(B => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b0 && CI1==1'b1 && CS==1'b1)
(B => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b0)
(B => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b1)
(B => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b0)
(B => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b1)
(B => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b1 && CI1==1'b0 && CS==1'b0)
(B => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b1 && CI1==1'b0 && CS==1'b1)
(B => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0==1'b0 && CS==1'b0)
(CI1 => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0==1'b0 && CS==1'b1)
(CI1 => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0==1'b1 && CS==1'b0)
(CI1 => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0==1'b1 && CS==1'b1)
(CI1 => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0==1'b0 && CS==1'b0)
(CI1 => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0==1'b0 && CS==1'b1)
(CI1 => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0==1'b1 && CS==1'b0)
(CI1 => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0==1'b1 && CS==1'b1)
(CI1 => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b0 && CI1==1'b1 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b0 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b1 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b1 && CI1==1'b0 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b0 && CI1==1'b0 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b0 && CI1==1'b0 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b0 && CI1==1'b1 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b0 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b1 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b1 && CI1==1'b0 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b1 && CI1==1'b1 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b1 && CI1==1'b1 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b0 && CI1==1'b1 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b0 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b1 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b1 && CI1==1'b0 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b0 && CI1==1'b0 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b0 && CI1==1'b0 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b0 && CI1==1'b1 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b0 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b1 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b1 && CI1==1'b0 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b1 && CI1==1'b1 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b1 && CI1==1'b1 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1==1'b0)
(CI0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1==1'b1)
(CI0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1==1'b0)
(CI0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1==1'b1)
(CI0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI1==1'b0)
(CI0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI1==1'b1)
(CI0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI1==1'b0)
(CI0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI1==1'b1)
(CI0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0==1'b0)
(CI1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0==1'b1)
(CI1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0==1'b0)
(CI1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0==1'b1)
(CI1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI0==1'b0)
(CI1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI0==1'b1)
(CI1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI0==1'b0)
(CI1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI0==1'b1)
(CI1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI0==1'b1 && CI1==1'b0)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0==1'b0 && CI1==1'b1)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0==1'b0 && CI1==1'b1)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI0==1'b1 && CI1==1'b0)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI0==1'b0 && CI1==1'b1)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0==1'b1 && CI1==1'b0)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0==1'b1 && CI1==1'b0)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI0==1'b0 && CI1==1'b1)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AFCSHCONX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AFCSHCONX4 (CO0N, CO1N, S, VDD, VSS, A, B, CI0, CI1, CS);
inout VDD, VSS;
output S, CO0N, CO1N;
input A, B, CI0, CI1, CS;
  xor I2 (s1, A, B, CI1);
  xor I3 (s2, A, B, CI0);
  and I4 (s3, CS, s1);
  not I5 (csn, CS);
  and I6 (s4, csn, s2);
  or I7 (sum_temp, s3, s4);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I8 (a_and_b, A, B);
  and I9 (a_and_ci0, A, CI0);
  and I10 (b_and_ci0, B, CI0);
  or I11 (cout0, a_and_b, a_and_ci0, b_and_ci0);
  and I12 (a_and_ci1, A, CI1);
  and I13 (b_and_ci1, B, CI1);
  or I14 (cout1, a_and_b, a_and_ci1, b_and_ci1);
  not I15 (cout0n_temp, cout0);
  assign CO0N = ((VDD === 1'b1) && (VSS === 1'b0))? cout0n_temp : 1'bx;
  not I16 (cout1n_temp, cout1);
  assign CO1N = ((VDD === 1'b1) && (VSS === 1'b0))? cout1n_temp : 1'bx;


specify
if (B==1'b0 && CI0==1'b1 && CI1==1'b0 && CS==1'b0)
(A => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b0 && CS==1'b1)
(A => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b0)
(A => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b1)
(A => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b0)
(A => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b1)
(A => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b1 && CS==1'b0)
(A => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b1 && CS==1'b1)
(A => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b0 && CS==1'b0)
(B => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b0 && CS==1'b1)
(B => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b0)
(B => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b1)
(B => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b0)
(B => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b1)
(B => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b1 && CS==1'b0)
(B => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b1 && CS==1'b1)
(B => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1==1'b0 && CS==1'b0)
(CI0 => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1==1'b0 && CS==1'b1)
(CI0 => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1==1'b1 && CS==1'b0)
(CI0 => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1==1'b1 && CS==1'b1)
(CI0 => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1==1'b0 && CS==1'b0)
(CI0 => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1==1'b0 && CS==1'b1)
(CI0 => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1==1'b1 && CS==1'b0)
(CI0 => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1==1'b1 && CS==1'b1)
(CI0 => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b0 && CI1==1'b1 && CS==1'b0)
(A => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b0 && CI1==1'b1 && CS==1'b1)
(A => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b0)
(A => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b1)
(A => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b0)
(A => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b1)
(A => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b1 && CI1==1'b0 && CS==1'b0)
(A => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b1 && CI1==1'b0 && CS==1'b1)
(A => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b0 && CI1==1'b1 && CS==1'b0)
(B => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b0 && CI1==1'b1 && CS==1'b1)
(B => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b0)
(B => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b1)
(B => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b0)
(B => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b1)
(B => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b1 && CI1==1'b0 && CS==1'b0)
(B => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b1 && CI1==1'b0 && CS==1'b1)
(B => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0==1'b0 && CS==1'b0)
(CI1 => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0==1'b0 && CS==1'b1)
(CI1 => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0==1'b1 && CS==1'b0)
(CI1 => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0==1'b1 && CS==1'b1)
(CI1 => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0==1'b0 && CS==1'b0)
(CI1 => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0==1'b0 && CS==1'b1)
(CI1 => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0==1'b1 && CS==1'b0)
(CI1 => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0==1'b1 && CS==1'b1)
(CI1 => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b0 && CI1==1'b1 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b0 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b1 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b1 && CI1==1'b0 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b0 && CI1==1'b0 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b0 && CI1==1'b0 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b0 && CI1==1'b1 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b0 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b1 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b1 && CI1==1'b0 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b1 && CI1==1'b1 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b1 && CI1==1'b1 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b0 && CI1==1'b1 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b0 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b1 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b1 && CI1==1'b0 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b0 && CI1==1'b0 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b0 && CI1==1'b0 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b0 && CI1==1'b1 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b0 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b1 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b1 && CI1==1'b0 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b1 && CI1==1'b1 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b1 && CI1==1'b1 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1==1'b0)
(CI0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1==1'b1)
(CI0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1==1'b0)
(CI0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1==1'b1)
(CI0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI1==1'b0)
(CI0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI1==1'b1)
(CI0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI1==1'b0)
(CI0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI1==1'b1)
(CI0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0==1'b0)
(CI1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0==1'b1)
(CI1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0==1'b0)
(CI1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0==1'b1)
(CI1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI0==1'b0)
(CI1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI0==1'b1)
(CI1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI0==1'b0)
(CI1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI0==1'b1)
(CI1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI0==1'b1 && CI1==1'b0)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0==1'b0 && CI1==1'b1)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0==1'b0 && CI1==1'b1)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI0==1'b1 && CI1==1'b0)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI0==1'b0 && CI1==1'b1)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0==1'b1 && CI1==1'b0)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0==1'b1 && CI1==1'b0)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI0==1'b0 && CI1==1'b1)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AFCSHCONX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AFHCINX2 (CO, S, VDD, VSS, A, B, CIN);
inout VDD, VSS;
output S, CO;
input A, B, CIN;
  not I0 (ci, CIN);
  xor I1 (sum_temp, A, B, ci);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I2 (a_and_b, A, B);
  and I3 (a_and_ci, A, ci);
  and I4 (b_and_ci, B, ci);
  or I5 (cout_temp, a_and_b, a_and_ci, b_and_ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
if (B==1'b0 && CIN==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CIN==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CIN==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CIN => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CIN => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CIN => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CIN => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AFHCINX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AFHCINX4 (CO, S, VDD, VSS, A, B, CIN);
inout VDD, VSS;
output S, CO;
input A, B, CIN;
  not I0 (ci, CIN);
  xor I1 (sum_temp, A, B, ci);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I2 (a_and_b, A, B);
  and I3 (a_and_ci, A, ci);
  and I4 (b_and_ci, B, ci);
  or I5 (cout_temp, a_and_b, a_and_ci, b_and_ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
if (B==1'b0 && CIN==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CIN==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CIN==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CIN => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CIN => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CIN => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CIN => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AFHCINX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AFHCONX2 (CON, S, VDD, VSS, A, B, CI);
inout VDD, VSS;
output S, CON;
input A, B, CI;
  xor I0 (sum_temp, A, B, CI);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I1 (a_and_b, A, B);
  and I2 (a_and_ci, A, CI);
  and I3 (b_and_ci, B, CI);
  or I4 (cout, a_and_b, a_and_ci, b_and_ci);
  not I5 (coutn_temp, cout);
  assign CON = ((VDD === 1'b1) && (VSS === 1'b0))? coutn_temp : 1'bx;


specify
if (B==1'b0 && CI==1'b1)
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AFHCONX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AFHCONX4 (CON, S, VDD, VSS, A, B, CI);
inout VDD, VSS;
output S, CON;
input A, B, CI;
  xor I0 (sum_temp, A, B, CI);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I1 (a_and_b, A, B);
  and I2 (a_and_ci, A, CI);
  and I3 (b_and_ci, B, CI);
  or I4 (cout, a_and_b, a_and_ci, b_and_ci);
  not I5 (coutn_temp, cout);
  assign CON = ((VDD === 1'b1) && (VSS === 1'b0))? coutn_temp : 1'bx;


specify
if (B==1'b0 && CI==1'b1)
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AFHCONX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AHHCINX2 (CO, S, VDD, VSS, A, CIN);
inout VDD, VSS;
output S, CO;
input A, CIN;
  not I0 (ci, CIN);
  xor I1 (sum_temp, A, ci);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I2 (cout_temp, A, ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CIN => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge CIN => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AHHCINX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AHHCINX4 (CO, S, VDD, VSS, A, CIN);
inout VDD, VSS;
output S, CO;
input A, CIN;
  not I0 (ci, CIN);
  xor I1 (sum_temp, A, ci);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I2 (cout_temp, A, ci);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CIN => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge CIN => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AHHCINX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AHHCONX2 (CON, S, VDD, VSS, A, CI);
inout VDD, VSS;
output S, CON;
input A, CI;
  xor I0 (sum_temp, A, CI);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and  I1 (cout, A, CI);
  not I2 (coutn_temp, cout);
  assign CON = ((VDD === 1'b1) && (VSS === 1'b0))? coutn_temp : 1'bx;


specify
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CI => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge CI => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AHHCONX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AHHCONX4 (CON, S, VDD, VSS, A, CI);
inout VDD, VSS;
output S, CON;
input A, CI;
  xor I0 (sum_temp, A, CI);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and  I1 (cout, A, CI);
  not I2 (coutn_temp, cout);
  assign CON = ((VDD === 1'b1) && (VSS === 1'b0))? coutn_temp : 1'bx;


specify
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CI => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge CI => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AHHCONX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2X1 (Y, VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2X2 (Y, VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2X4 (Y, VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2XL (Y, VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  and (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3X1 (Y, VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  and (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3X2 (Y, VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  and (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3X4 (Y, VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  and (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3XL (Y, VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  and (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4X1 (Y, VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  and (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4X2 (Y, VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  and (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4X4 (Y, VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  and (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4XL (Y, VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  and (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ANTENNA (VDD, VSS, A);
 inout VDD, VSS;
input A;

specify

endspecify
endmodule // ANTENNA
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211X1 (Y, VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI211X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211X2 (Y, VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI211X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211X4 (Y, VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI211X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211XL (Y, VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI211XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21X1 (Y, VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21X2 (Y, VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21X4 (Y, VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21XL (Y, VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221X1 (Y, VDD, VSS, A0, A1, B0, B1, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(out_temp, C0, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI221X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221X2 (Y, VDD, VSS, A0, A1, B0, B1, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(out_temp, C0, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI221X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221X4 (Y, VDD, VSS, A0, A1, B0, B1, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(out_temp, C0, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI221X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221XL (Y, VDD, VSS, A0, A1, B0, B1, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(out_temp, C0, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI221XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222X1 (Y, VDD, VSS, A0, A1, B0, B1, C0, C1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(out_temp, outA, outB, outC);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI222X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222X2 (Y, VDD, VSS, A0, A1, B0, B1, C0, C1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(out_temp, outA, outB, outC);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI222X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222X4 (Y, VDD, VSS, A0, A1, B0, B1, C0, C1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(out_temp, outA, outB, outC);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI222X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222XL (Y, VDD, VSS, A0, A1, B0, B1, C0, C1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(out_temp, outA, outB, outC);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI222XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22X1 (Y, VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22X2 (Y, VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22X4 (Y, VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22XL (Y, VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB1X1 (Y, VDD, VSS, A0N, A1N, B0);
inout VDD, VSS;
output Y;
input A0N, A1N, B0;



  nor I0 (outA, A0N, A1N);
  nor I1 (out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB1X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB1X2 (Y, VDD, VSS, A0N, A1N, B0);
inout VDD, VSS;
output Y;
input A0N, A1N, B0;



  nor I0 (outA, A0N, A1N);
  nor I1 (out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB1X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB1X4 (Y, VDD, VSS, A0N, A1N, B0);
inout VDD, VSS;
output Y;
input A0N, A1N, B0;



  nor I0 (outA, A0N, A1N);
  nor I1 (out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB1X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB1XL (Y, VDD, VSS, A0N, A1N, B0);
inout VDD, VSS;
output Y;
input A0N, A1N, B0;



  nor I0 (outA, A0N, A1N);
  nor I1 (out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB1XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB2X1 (Y, VDD, VSS, A0N, A1N, B0, B1);
inout VDD, VSS;
output Y;
input A0N, A1N, B0, B1;



  nor I0 (outA, A0N, A1N);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB2X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB2X2 (Y, VDD, VSS, A0N, A1N, B0, B1);
inout VDD, VSS;
output Y;
input A0N, A1N, B0, B1;



  nor I0 (outA, A0N, A1N);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB2X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB2X4 (Y, VDD, VSS, A0N, A1N, B0, B1);
inout VDD, VSS;
output Y;
input A0N, A1N, B0, B1;



  nor I0 (outA, A0N, A1N);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB2X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB2XL (Y, VDD, VSS, A0N, A1N, B0, B1);
inout VDD, VSS;
output Y;
input A0N, A1N, B0, B1;



  nor I0 (outA, A0N, A1N);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB2XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31X1 (Y, VDD, VSS, A0, A1, A2, B0);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI31X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31X2 (Y, VDD, VSS, A0, A1, A2, B0);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI31X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31X4 (Y, VDD, VSS, A0, A1, A2, B0);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI31X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31XL (Y, VDD, VSS, A0, A1, A2, B0);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI31XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32X1 (Y, VDD, VSS, A0, A1, A2, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI32X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32X2 (Y, VDD, VSS, A0, A1, A2, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI32X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32X4 (Y, VDD, VSS, A0, A1, A2, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI32X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32XL (Y, VDD, VSS, A0, A1, A2, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI32XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI33X1 (Y, VDD, VSS, A0, A1, A2, B0, B1, B2);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1, B2;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1, B2);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI33X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI33X2 (Y, VDD, VSS, A0, A1, A2, B0, B1, B2);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1, B2;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1, B2);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI33X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI33X4 (Y, VDD, VSS, A0, A1, A2, B0, B1, B2);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1, B2;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1, B2);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI33X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI33XL (Y, VDD, VSS, A0, A1, A2, B0, B1, B2);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1, B2;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1, B2);
  nor I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI33XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BENCX1 (A, S, X2, VDD, VSS, M0, M1, M2);
inout VDD, VSS;
output S, A, X2;
input M2, M1, M0;

  not I0 (m1n, M1);
  not I1 (m0n, M0);
  or  I3 (m1n_or_m0n, m1n, m0n);
  nand I4 (subb_temp, M2, m1n_or_m0n);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? subb_temp : 1'bx;
  or  I5 (m1_or_m0, M1, M0);
  nand I6 (addb_temp, m2n, m1_or_m0);
  assign A = ((VDD === 1'b1) && (VSS === 1'b0))? addb_temp : 1'bx;
  xor I7 (x2n, M1, M0);
  not I8 (x2_temp, x2n);
  assign X2 = ((VDD === 1'b1) && (VSS === 1'b0))? x2_temp : 1'bx;
  not I9 (m2n, M2);



specify
(M0 => A) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => A) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => A) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => A) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b1)
(M2 => A) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b0)
(M2 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BENCX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BENCX2 (A, S, X2, VDD, VSS, M0, M1, M2);
inout VDD, VSS;
output S, A, X2;
input M2, M1, M0;

  not I0 (m1n, M1);
  not I1 (m0n, M0);
  or  I3 (m1n_or_m0n, m1n, m0n);
  nand I4 (subb_temp, M2, m1n_or_m0n);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? subb_temp : 1'bx;
  or  I5 (m1_or_m0, M1, M0);
  nand I6 (addb_temp, m2n, m1_or_m0);
  assign A = ((VDD === 1'b1) && (VSS === 1'b0))? addb_temp : 1'bx;
  xor I7 (x2n, M1, M0);
  not I8 (x2_temp, x2n);
  assign X2 = ((VDD === 1'b1) && (VSS === 1'b0))? x2_temp : 1'bx;
  not I9 (m2n, M2);



specify
(M0 => A) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => A) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => A) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => A) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b1)
(M2 => A) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b0)
(M2 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BENCX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BENCX4 (A, S, X2, VDD, VSS, M0, M1, M2);
inout VDD, VSS;
output S, A, X2;
input M2, M1, M0;

  not I0 (m1n, M1);
  not I1 (m0n, M0);
  or  I3 (m1n_or_m0n, m1n, m0n);
  nand I4 (subb_temp, M2, m1n_or_m0n);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? subb_temp : 1'bx;
  or  I5 (m1_or_m0, M1, M0);
  nand I6 (addb_temp, m2n, m1_or_m0);
  assign A = ((VDD === 1'b1) && (VSS === 1'b0))? addb_temp : 1'bx;
  xor I7 (x2n, M1, M0);
  not I8 (x2_temp, x2n);
  assign X2 = ((VDD === 1'b1) && (VSS === 1'b0))? x2_temp : 1'bx;
  not I9 (m2n, M2);



specify
(M0 => A) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => A) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => A) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => A) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b1)
(M2 => A) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b0)
(M2 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BENCX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BMXX1 (PP, VDD, VSS, A, M0, M1, S, X2);
inout VDD, VSS;
output PP;
input X2, A, S, M1, M0;

  udp_bmx I0 (z_temp, X2, A, S, M1, M0);
  assign PP = ((VDD === 1'b1) && (VSS === 1'b0))? z_temp : 1'bx;



specify
if (M0==1'b0 && M1==1'b1 && S==1'b0 && X2==1'b0)
(A => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1 && S==1'b1 && X2==1'b0)
(A => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0 && S==1'b0 && X2==1'b1)
(A => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0 && S==1'b1 && X2==1'b1)
(A => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b1 && S==1'b0 && X2==1'b0)
(A => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b1 && S==1'b0 && X2==1'b1)
(A => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b1 && S==1'b1 && X2==1'b0)
(A => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b1 && S==1'b1 && X2==1'b1)
(A => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M1==1'b0)
(posedge M0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M1==1'b0)
(negedge M0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M1==1'b1)
(posedge M0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M1==1'b1)
(negedge M0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0)
(posedge M1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0)
(negedge M1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1)
(posedge M1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1)
(negedge M1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && M0==1'b0 && M1==1'b0 && X2==1'b0)
(S => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && M0==1'b0 && M1==1'b0 && X2==1'b1)
(S => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && M0==1'b0 && M1==1'b1 && X2==1'b1)
(S => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && M0==1'b1 && M1==1'b0 && X2==1'b0)
(S => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && M0==1'b0 && M1==1'b0 && X2==1'b0)
(S => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && M0==1'b0 && M1==1'b0 && X2==1'b1)
(S => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && M0==1'b0 && M1==1'b1 && X2==1'b1)
(S => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && M0==1'b1 && M1==1'b0 && X2==1'b0)
(S => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && M0==1'b0 && M1==1'b1 && S==1'b1)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && M0==1'b1 && M1==1'b0 && S==1'b0)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && M0==1'b1 && M1==1'b0 && S==1'b1)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && M0==1'b0 && M1==1'b1 && S==1'b0)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BMXX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFX1 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFX12 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFX12
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFX16 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFX16
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFX2 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFX20 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFX20
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFX3 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFX3
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFX4 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFX8 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFX8
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFXL (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUFX1 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUFX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUFX12 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUFX12
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUFX16 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUFX16
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUFX2 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUFX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUFX20 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUFX20
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUFX3 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUFX3
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUFX4 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUFX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUFX8 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUFX8
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUFXL (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUFXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINVX1 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINVX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINVX12 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINVX12
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINVX16 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINVX16
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINVX2 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINVX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINVX20 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINVX20
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINVX3 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINVX3
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINVX4 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINVX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINVX8 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINVX8
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINVXL (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINVXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CMPR22X1 (CO, S, VDD, VSS, A, B);
inout VDD, VSS;
output S, CO;
input A, B;
  xor I0(sum_temp, A, B);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I1(cout_temp, A, B);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;


specify
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CMPR22X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CMPR32X1 (CO, S, VDD, VSS, A, B, C);
inout VDD, VSS;
output S, CO;
input A, B, C;

  xor I0 (t1, A, B);
  xor I1 (sum_temp, t1, C);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? sum_temp : 1'bx;
  and I2 (t2, A, B);
  and I3 (t3, t1, C);
  or  I4 (cout_temp, t2, t3);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? cout_temp : 1'bx;



specify
if (B==1'b0 && C==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CMPR32X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CMPR42X1 (CO, ICO, S, VDD, VSS, A, B, C, D, ICI);
inout VDD, VSS;
output S, CO, ICO;
input A, B, C, D, ICI;

  xor I0 (t1, A, B);
  xor I1 (IS, t1, C);
  and I2 (t2, A, B);
  and I3 (t3, A, C);
  and I4 (t4, B, C);
  or   I5 (co_temp, t2, t3, t4);
  assign ICO = ((VDD === 1'b1) && (VSS === 1'b0))? co_temp : 1'bx;
  xor I6 (ss, IS, D);
  xor  I7 (S_temp, ss, ICI);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? S_temp : 1'bx;
  and I8 (t5, IS, D);
  and I9 (t6, IS, ICI);
  and I10 (t7, D, ICI);
  or   I11 (c_temp, t5, t6, t7);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? c_temp : 1'bx;



specify
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0 && ICI==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1 && ICI==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0 && ICI==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1 && ICI==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && ICI==1'b1)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && ICI==1'b0)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && ICI==1'b0)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && ICI==1'b1)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && ICI==1'b0)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && ICI==1'b1)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && ICI==1'b1)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && ICI==1'b0)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && ICI==1'b0)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && ICI==1'b1)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && ICI==1'b1)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && ICI==1'b0)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && ICI==1'b1)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && ICI==1'b0)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && ICI==1'b0)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && ICI==1'b1)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b0)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b1)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CMPR42X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CMPR42X2 (CO, ICO, S, VDD, VSS, A, B, C, D, ICI);
inout VDD, VSS;
output S, CO, ICO;
input A, B, C, D, ICI;

  xor I0 (t1, A, B);
  xor I1 (IS, t1, C);
  and I2 (t2, A, B);
  and I3 (t3, A, C);
  and I4 (t4, B, C);
  or   I5 (co_temp, t2, t3, t4);
  assign ICO = ((VDD === 1'b1) && (VSS === 1'b0))? co_temp : 1'bx;
  xor I6 (ss, IS, D);
  xor  I7 (S_temp, ss, ICI);
  assign S = ((VDD === 1'b1) && (VSS === 1'b0))? S_temp : 1'bx;
  and I8 (t5, IS, D);
  and I9 (t6, IS, ICI);
  and I10 (t7, D, ICI);
  or   I11 (c_temp, t5, t6, t7);
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0))? c_temp : 1'bx;



specify
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0 && ICI==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1 && ICI==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0 && ICI==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1 && ICI==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && ICI==1'b1)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && ICI==1'b0)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && ICI==1'b0)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && ICI==1'b1)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && ICI==1'b0)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && ICI==1'b1)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && ICI==1'b1)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && ICI==1'b0)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && ICI==1'b0)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && ICI==1'b1)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && ICI==1'b1)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && ICI==1'b0)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && ICI==1'b1)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && ICI==1'b0)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && ICI==1'b0)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && ICI==1'b1)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b0)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b1)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CMPR42X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DFFHQX1 (Q, VDD, VSS, CK, D);
inout VDD, VSS;
output Q;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);


specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFHQX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFHQX2 (Q, VDD, VSS, CK, D);
inout VDD, VSS;
output Q;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);


specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFHQX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFHQX4 (Q, VDD, VSS, CK, D);
inout VDD, VSS;
output Q;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);


specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFHQX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFHQXL (Q, VDD, VSS, CK, D);
inout VDD, VSS;
output Q;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);


specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFHQXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNRX1 (Q, QN, VDD, VSS, CKN, D, RN);
inout VDD, VSS;
output Q, QN;
input  D, CKN, RN;
reg NOTIFIER;
supply1 xSN;

  buf   XX0 (xRN, RN);
  not      IC (clk, CKN);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_D ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, negedge CKN &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // DFFNRX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNRX2 (Q, QN, VDD, VSS, CKN, D, RN);
inout VDD, VSS;
output Q, QN;
input  D, CKN, RN;
reg NOTIFIER;
supply1 xSN;

  buf   XX0 (xRN, RN);
  not      IC (clk, CKN);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_D ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, negedge CKN &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // DFFNRX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNRX4 (Q, QN, VDD, VSS, CKN, D, RN);
inout VDD, VSS;
output Q, QN;
input  D, CKN, RN;
reg NOTIFIER;
supply1 xSN;

  buf   XX0 (xRN, RN);
  not      IC (clk, CKN);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_D ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, negedge CKN &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // DFFNRX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNRXL (Q, QN, VDD, VSS, CKN, D, RN);
inout VDD, VSS;
output Q, QN;
input  D, CKN, RN;
reg NOTIFIER;
supply1 xSN;

  buf   XX0 (xRN, RN);
  not      IC (clk, CKN);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_D ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, negedge CKN &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // DFFNRXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSRX1 (Q, QN, VDD, VSS, CKN, D, RN, SN);
inout VDD, VSS;
output Q, QN;
input  D, CKN, SN, RN;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  not      IC (clk, CKN);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, negedge CKN &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFNSRX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSRX2 (Q, QN, VDD, VSS, CKN, D, RN, SN);
inout VDD, VSS;
output Q, QN;
input  D, CKN, SN, RN;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  not      IC (clk, CKN);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, negedge CKN &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFNSRX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSRX4 (Q, QN, VDD, VSS, CKN, D, RN, SN);
inout VDD, VSS;
output Q, QN;
input  D, CKN, SN, RN;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  not      IC (clk, CKN);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, negedge CKN &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFNSRX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSRXL (Q, QN, VDD, VSS, CKN, D, RN, SN);
inout VDD, VSS;
output Q, QN;
input  D, CKN, SN, RN;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  not      IC (clk, CKN);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, negedge CKN &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFNSRXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSX1 (Q, QN, VDD, VSS, CKN, D, SN);
inout VDD, VSS;
output Q, QN;
input  D, CKN, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  not      IC (clk, CKN);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFNSX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSX2 (Q, QN, VDD, VSS, CKN, D, SN);
inout VDD, VSS;
output Q, QN;
input  D, CKN, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  not      IC (clk, CKN);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFNSX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSX4 (Q, QN, VDD, VSS, CKN, D, SN);
inout VDD, VSS;
output Q, QN;
input  D, CKN, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  not      IC (clk, CKN);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFNSX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSXL (Q, QN, VDD, VSS, CKN, D, SN);
inout VDD, VSS;
output Q, QN;
input  D, CKN, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  not      IC (clk, CKN);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFNSXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNX1 (Q, QN, VDD, VSS, CKN, D);
inout VDD, VSS;
output Q, QN;
input  D, CKN;
reg NOTIFIER;
supply1 xSN,xRN;
  not      IC (clk, CKN);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);


specify
$width(posedge CKN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFNX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNX2 (Q, QN, VDD, VSS, CKN, D);
inout VDD, VSS;
output Q, QN;
input  D, CKN;
reg NOTIFIER;
supply1 xSN,xRN;
  not      IC (clk, CKN);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);


specify
$width(posedge CKN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFNX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNX4 (Q, QN, VDD, VSS, CKN, D);
inout VDD, VSS;
output Q, QN;
input  D, CKN;
reg NOTIFIER;
supply1 xSN,xRN;
  not      IC (clk, CKN);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);


specify
$width(posedge CKN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFNX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNXL (Q, QN, VDD, VSS, CKN, D);
inout VDD, VSS;
output Q, QN;
input  D, CKN;
reg NOTIFIER;
supply1 xSN,xRN;
  not      IC (clk, CKN);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);


specify
$width(posedge CKN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFNXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRHQX1 (Q, VDD, VSS, CK, D, RN);
inout VDD, VSS;
output Q;
input  D, CK, RN;
reg NOTIFIER;
supply1 xSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_RN ;
wire ENABLE_D ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFRHQX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRHQX2 (Q, VDD, VSS, CK, D, RN);
inout VDD, VSS;
output Q;
input  D, CK, RN;
reg NOTIFIER;
supply1 xSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_RN ;
wire ENABLE_D ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFRHQX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRHQX4 (Q, VDD, VSS, CK, D, RN);
inout VDD, VSS;
output Q;
input  D, CK, RN;
reg NOTIFIER;
supply1 xSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_RN ;
wire ENABLE_D ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFRHQX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRHQXL (Q, VDD, VSS, CK, D, RN);
inout VDD, VSS;
output Q;
input  D, CK, RN;
reg NOTIFIER;
supply1 xSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_RN ;
wire ENABLE_D ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFRHQXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRX1 (Q, QN, VDD, VSS, CK, D, RN);
inout VDD, VSS;
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
supply1 xSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_D ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // DFFRX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRX2 (Q, QN, VDD, VSS, CK, D, RN);
inout VDD, VSS;
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
supply1 xSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_D ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // DFFRX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRX4 (Q, QN, VDD, VSS, CK, D, RN);
inout VDD, VSS;
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
supply1 xSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_D ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // DFFRX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRXL (Q, QN, VDD, VSS, CK, D, RN);
inout VDD, VSS;
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
supply1 xSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_D ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // DFFRXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSHQX1 (Q, VDD, VSS, CK, D, SN);
inout VDD, VSS;
output Q;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // DFFSHQX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSHQX2 (Q, VDD, VSS, CK, D, SN);
inout VDD, VSS;
output Q;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // DFFSHQX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSHQX4 (Q, VDD, VSS, CK, D, SN);
inout VDD, VSS;
output Q;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // DFFSHQX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSHQXL (Q, VDD, VSS, CK, D, SN);
inout VDD, VSS;
output Q;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // DFFSHQXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRHQX1 (Q, VDD, VSS, CK, D, RN, SN);
inout VDD, VSS;
output Q;
input  D, CK, SN, RN;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // DFFSRHQX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRHQX2 (Q, VDD, VSS, CK, D, RN, SN);
inout VDD, VSS;
output Q;
input  D, CK, SN, RN;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // DFFSRHQX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRHQX4 (Q, VDD, VSS, CK, D, RN, SN);
inout VDD, VSS;
output Q;
input  D, CK, SN, RN;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // DFFSRHQX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRHQXL (Q, VDD, VSS, CK, D, RN, SN);
inout VDD, VSS;
output Q;
input  D, CK, SN, RN;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // DFFSRHQXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRX1 (Q, QN, VDD, VSS, CK, D, RN, SN);
inout VDD, VSS;
output Q, QN;
input  D, CK, SN, RN;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSRX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRX2 (Q, QN, VDD, VSS, CK, D, RN, SN);
inout VDD, VSS;
output Q, QN;
input  D, CK, SN, RN;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSRX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRX4 (Q, QN, VDD, VSS, CK, D, RN, SN);
inout VDD, VSS;
output Q, QN;
input  D, CK, SN, RN;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSRX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRXL (Q, QN, VDD, VSS, CK, D, RN, SN);
inout VDD, VSS;
output Q, QN;
input  D, CK, SN, RN;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSRXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSX1 (Q, QN, VDD, VSS, CK, D, SN);
inout VDD, VSS;
output Q, QN;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSX2 (Q, QN, VDD, VSS, CK, D, SN);
inout VDD, VSS;
output Q, QN;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSX4 (Q, QN, VDD, VSS, CK, D, SN);
inout VDD, VSS;
output Q, QN;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSXL (Q, QN, VDD, VSS, CK, D, SN);
inout VDD, VSS;
output Q, QN;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFTRX1 (Q, QN, VDD, VSS, CK, D, RN);
inout VDD, VSS;
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
supply1 xSN, EN,flag;

  buf   XX0 (xRN, RN);
  and F0 (rn_and_sn, xRN,xSN);
  buf     IC (clk, CK);
  udp_edfft_PWR  I0 (n0, D, clk, xRN, xSN, EN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_D ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (RN==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (RN==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFTRX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFTRX2 (Q, QN, VDD, VSS, CK, D, RN);
inout VDD, VSS;
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
supply1 xSN, EN,flag;

  buf   XX0 (xRN, RN);
  and F0 (rn_and_sn, xRN,xSN);
  buf     IC (clk, CK);
  udp_edfft_PWR  I0 (n0, D, clk, xRN, xSN, EN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_D ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (RN==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (RN==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFTRX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFTRX4 (Q, QN, VDD, VSS, CK, D, RN);
inout VDD, VSS;
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
supply1 xSN, EN,flag;

  buf   XX0 (xRN, RN);
  and F0 (rn_and_sn, xRN,xSN);
  buf     IC (clk, CK);
  udp_edfft_PWR  I0 (n0, D, clk, xRN, xSN, EN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_D ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (RN==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (RN==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFTRX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFTRXL (Q, QN, VDD, VSS, CK, D, RN);
inout VDD, VSS;
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
supply1 xSN, EN,flag;

  buf   XX0 (xRN, RN);
  and F0 (rn_and_sn, xRN,xSN);
  buf     IC (clk, CK);
  udp_edfft_PWR  I0 (n0, D, clk, xRN, xSN, EN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_D ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (RN==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (RN==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFTRXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFX1 (Q, QN, VDD, VSS, CK, D);
inout VDD, VSS;
output Q, QN;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);


specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFX2 (Q, QN, VDD, VSS, CK, D);
inout VDD, VSS;
output Q, QN;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);


specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFX4 (Q, QN, VDD, VSS, CK, D);
inout VDD, VSS;
output Q, QN;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);


specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFXL (Q, QN, VDD, VSS, CK, D);
inout VDD, VSS;
output Q, QN;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);


specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DLY1X1 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLY1X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLY2X1 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLY2X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLY3X1 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLY3X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLY4X1 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  buf I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLY4X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module EDFFTRX1 (Q, QN, VDD, VSS, CK, D, E, RN);
inout VDD, VSS;
output Q, QN;
input D, CK, E, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

  udp_edfft_PWR  I0 (n0, D, CK, xRN, xSN, E, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_E_OR_NOT_RN ;
wire ENABLE_E_AND_RN ;
wire ENABLE_RN ;
wire ENABLE_D_OR_NOT_E ;
assign ENABLE_E_OR_NOT_RN = (E | !RN) ? 1'b1:1'b0;
assign ENABLE_E_AND_RN = (E&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D_OR_NOT_E = (D | !E) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_NOT_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_NOT_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_OR_NOT_E == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_OR_NOT_E == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (E==1'b1 && RN==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFFTRX1
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFFTRX2 (Q, QN, VDD, VSS, CK, D, E, RN);
inout VDD, VSS;
output Q, QN;
input D, CK, E, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

  udp_edfft_PWR  I0 (n0, D, CK, xRN, xSN, E, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_E_OR_NOT_RN ;
wire ENABLE_E_AND_RN ;
wire ENABLE_RN ;
wire ENABLE_D_OR_NOT_E ;
assign ENABLE_E_OR_NOT_RN = (E | !RN) ? 1'b1:1'b0;
assign ENABLE_E_AND_RN = (E&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D_OR_NOT_E = (D | !E) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_NOT_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_NOT_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_OR_NOT_E == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_OR_NOT_E == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (E==1'b1 && RN==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFFTRX2
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFFTRX4 (Q, QN, VDD, VSS, CK, D, E, RN);
inout VDD, VSS;
output Q, QN;
input D, CK, E, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

  udp_edfft_PWR  I0 (n0, D, CK, xRN, xSN, E, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_E_OR_NOT_RN ;
wire ENABLE_E_AND_RN ;
wire ENABLE_RN ;
wire ENABLE_D_OR_NOT_E ;
assign ENABLE_E_OR_NOT_RN = (E | !RN) ? 1'b1:1'b0;
assign ENABLE_E_AND_RN = (E&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D_OR_NOT_E = (D | !E) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_NOT_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_NOT_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_OR_NOT_E == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_OR_NOT_E == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (E==1'b1 && RN==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFFTRX4
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFFTRXL (Q, QN, VDD, VSS, CK, D, E, RN);
inout VDD, VSS;
output Q, QN;
input D, CK, E, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

  udp_edfft_PWR  I0 (n0, D, CK, xRN, xSN, E, VDD, VSS, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_E_OR_NOT_RN ;
wire ENABLE_E_AND_RN ;
wire ENABLE_RN ;
wire ENABLE_D_OR_NOT_E ;
assign ENABLE_E_OR_NOT_RN = (E | !RN) ? 1'b1:1'b0;
assign ENABLE_E_AND_RN = (E&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D_OR_NOT_E = (D | !E) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_NOT_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_NOT_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_OR_NOT_E == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_OR_NOT_E == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (E==1'b1 && RN==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFFTRXL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFFX1 (Q, QN, VDD, VSS, CK, D, E);
inout VDD, VSS;
output Q, QN;
input D, CK, E;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff_PWR  I0 (n0, D, CK, xRN, xSN, E, VDD, VSS, NOTIFIER);
  buf     B1 (Q, n0);
  not      I1 (QN, n0);

wire ENABLE_E ;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFFX1
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFFX2 (Q, QN, VDD, VSS, CK, D, E);
inout VDD, VSS;
output Q, QN;
input D, CK, E;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff_PWR  I0 (n0, D, CK, xRN, xSN, E, VDD, VSS, NOTIFIER);
  buf     B1 (Q, n0);
  not      I1 (QN, n0);

wire ENABLE_E ;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFFX2
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFFX4 (Q, QN, VDD, VSS, CK, D, E);
inout VDD, VSS;
output Q, QN;
input D, CK, E;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff_PWR  I0 (n0, D, CK, xRN, xSN, E, VDD, VSS, NOTIFIER);
  buf     B1 (Q, n0);
  not      I1 (QN, n0);

wire ENABLE_E ;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFFX4
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFFXL (Q, QN, VDD, VSS, CK, D, E);
inout VDD, VSS;
output Q, QN;
input D, CK, E;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff_PWR  I0 (n0, D, CK, xRN, xSN, E, VDD, VSS, NOTIFIER);
  buf     B1 (Q, n0);
  not      I1 (QN, n0);

wire ENABLE_E ;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFFXL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module FILL1 (VDD, VSS);
inout VDD, VSS;
endmodule //FILL1

`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILL16 (VDD, VSS);
inout VDD, VSS;
endmodule //FILL16

`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILL2 (VDD, VSS);
inout VDD, VSS;
endmodule //FILL2

`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILL32 (VDD, VSS);
inout VDD, VSS;
endmodule //FILL32

`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILL4 (VDD, VSS);
inout VDD, VSS;
endmodule //FILL4

`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILL64 (VDD, VSS);
inout VDD, VSS;
endmodule //FILL64

`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILL8 (VDD, VSS);
inout VDD, VSS;
endmodule //FILL8

`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILLCAP16 (VDD, VSS);
inout VDD, VSS;

specify

endspecify
endmodule // FILLCAP16
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILLCAP3 (VDD, VSS);
inout VDD, VSS;

specify

endspecify
endmodule // FILLCAP3
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILLCAP32 (VDD, VSS);
inout VDD, VSS;

specify

endspecify
endmodule // FILLCAP32
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILLCAP4 (VDD, VSS);
inout VDD, VSS;

specify

endspecify
endmodule // FILLCAP4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILLCAP5 (VDD, VSS);
inout VDD, VSS;

specify

endspecify
endmodule // FILLCAP5
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILLCAP64 (VDD, VSS);
inout VDD, VSS;

specify

endspecify
endmodule // FILLCAP64
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILLCAP8 (VDD, VSS);
inout VDD, VSS;

specify

endspecify
endmodule // FILLCAP8
`endcelldefine
`timescale 1ns/1ps
`celldefine
module HOLDX1 (VDD, VSS, Y);
inout VDD, VSS;
inout Y;

wire io_wire;

  assign io_wire = ((VDD === 1'b1) && (VSS === 1'b0))? Y : 1'bx;
  buf(weak0,weak1) I0(Y, io_wire);



specify

endspecify
endmodule // HOLDX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INVX1 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INVX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INVX12 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INVX12
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INVX16 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INVX16
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INVX2 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INVX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INVX20 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INVX20
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INVX3 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INVX3
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INVX4 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INVX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INVX8 (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INVX8
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INVXL (Y, VDD, VSS, A);
inout VDD, VSS;
output Y;
input A;

  not I0(out_temp, A);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INVXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module JKFFRX1 (Q, QN, VDD, VSS, CK, J, K, RN);
inout VDD, VSS;
output Q, QN;
input  J, K, CK, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);

udp_jkff_PWR  I0 (n0,J, K,CK,xRN,xSN,VDD, VSS, NOTIFIER); 
buf I1 (Q,n0);
not I2 (QN,n0);

wire ENABLE_J_AND_RN_OR_K_AND_RN ;
wire ENABLE_RN ;
wire ENABLE_J ;
assign ENABLE_J_AND_RN_OR_K_AND_RN = (J&RN | K&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_J = (J) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_J_AND_RN_OR_K_AND_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_J_AND_RN_OR_K_AND_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_J == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // JKFFRX1
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFRX2 (Q, QN, VDD, VSS, CK, J, K, RN);
inout VDD, VSS;
output Q, QN;
input  J, K, CK, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);

udp_jkff_PWR  I0 (n0,J, K,CK,xRN,xSN,VDD, VSS, NOTIFIER); 
buf I1 (Q,n0);
not I2 (QN,n0);

wire ENABLE_J_AND_RN_OR_K_AND_RN ;
wire ENABLE_RN ;
wire ENABLE_J ;
assign ENABLE_J_AND_RN_OR_K_AND_RN = (J&RN | K&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_J = (J) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_J_AND_RN_OR_K_AND_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_J_AND_RN_OR_K_AND_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_J == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // JKFFRX2
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFRX4 (Q, QN, VDD, VSS, CK, J, K, RN);
inout VDD, VSS;
output Q, QN;
input  J, K, CK, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);

udp_jkff_PWR  I0 (n0,J, K,CK,xRN,xSN,VDD, VSS, NOTIFIER); 
buf I1 (Q,n0);
not I2 (QN,n0);

wire ENABLE_J_AND_RN_OR_K_AND_RN ;
wire ENABLE_RN ;
wire ENABLE_J ;
assign ENABLE_J_AND_RN_OR_K_AND_RN = (J&RN | K&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_J = (J) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_J_AND_RN_OR_K_AND_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_J_AND_RN_OR_K_AND_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_J == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // JKFFRX4
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFRXL (Q, QN, VDD, VSS, CK, J, K, RN);
inout VDD, VSS;
output Q, QN;
input  J, K, CK, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);

udp_jkff_PWR  I0 (n0,J, K,CK,xRN,xSN,VDD, VSS, NOTIFIER); 
buf I1 (Q,n0);
not I2 (QN,n0);

wire ENABLE_J_AND_RN_OR_K_AND_RN ;
wire ENABLE_RN ;
wire ENABLE_J ;
assign ENABLE_J_AND_RN_OR_K_AND_RN = (J&RN | K&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_J = (J) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_J_AND_RN_OR_K_AND_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_J_AND_RN_OR_K_AND_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_J == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // JKFFRXL
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFSRX1 (Q, QN, VDD, VSS, CK, J, K, RN, SN);
inout VDD, VSS;
output Q, QN;
input  J, K, CK, SN, RN;
reg NOTIFIER;

  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);

udp_jkff_PWR  I0 (n0,J, K,CK,xRN,xSN,VDD, VSS, NOTIFIER); 
buf I1 (Q,n0);
not I2 (QN,n0);

wire ENABLE_J_AND_RN_AND_SN_OR_K_AND_RN_AND_SN ;
wire ENABLE_RN_AND_SN ;
wire ENABLE_J_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_K_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_J_AND_RN_AND_SN_OR_K_AND_RN_AND_SN = (J&RN&SN | K&RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_J_AND_SN = (J&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_K_AND_RN = (K&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_J_AND_RN_AND_SN_OR_K_AND_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_J_AND_RN_AND_SN_OR_K_AND_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_J_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_K_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // JKFFSRX1
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFSRX2 (Q, QN, VDD, VSS, CK, J, K, RN, SN);
inout VDD, VSS;
output Q, QN;
input  J, K, CK, SN, RN;
reg NOTIFIER;

  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);

udp_jkff_PWR  I0 (n0,J, K,CK,xRN,xSN,VDD, VSS, NOTIFIER); 
buf I1 (Q,n0);
not I2 (QN,n0);

wire ENABLE_J_AND_RN_AND_SN_OR_K_AND_RN_AND_SN ;
wire ENABLE_RN_AND_SN ;
wire ENABLE_J_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_K_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_J_AND_RN_AND_SN_OR_K_AND_RN_AND_SN = (J&RN&SN | K&RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_J_AND_SN = (J&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_K_AND_RN = (K&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_J_AND_RN_AND_SN_OR_K_AND_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_J_AND_RN_AND_SN_OR_K_AND_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_J_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_K_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // JKFFSRX2
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFSRX4 (Q, QN, VDD, VSS, CK, J, K, RN, SN);
inout VDD, VSS;
output Q, QN;
input  J, K, CK, SN, RN;
reg NOTIFIER;

  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);

udp_jkff_PWR  I0 (n0,J, K,CK,xRN,xSN,VDD, VSS, NOTIFIER); 
buf I1 (Q,n0);
not I2 (QN,n0);

wire ENABLE_J_AND_RN_AND_SN_OR_K_AND_RN_AND_SN ;
wire ENABLE_RN_AND_SN ;
wire ENABLE_J_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_K_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_J_AND_RN_AND_SN_OR_K_AND_RN_AND_SN = (J&RN&SN | K&RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_J_AND_SN = (J&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_K_AND_RN = (K&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_J_AND_RN_AND_SN_OR_K_AND_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_J_AND_RN_AND_SN_OR_K_AND_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_J_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_K_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // JKFFSRX4
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFSRXL (Q, QN, VDD, VSS, CK, J, K, RN, SN);
inout VDD, VSS;
output Q, QN;
input  J, K, CK, SN, RN;
reg NOTIFIER;

  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);

udp_jkff_PWR  I0 (n0,J, K,CK,xRN,xSN,VDD, VSS, NOTIFIER); 
buf I1 (Q,n0);
not I2 (QN,n0);

wire ENABLE_J_AND_RN_AND_SN_OR_K_AND_RN_AND_SN ;
wire ENABLE_RN_AND_SN ;
wire ENABLE_J_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_K_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_J_AND_RN_AND_SN_OR_K_AND_RN_AND_SN = (J&RN&SN | K&RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_J_AND_SN = (J&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_K_AND_RN = (K&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_J_AND_RN_AND_SN_OR_K_AND_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_J_AND_RN_AND_SN_OR_K_AND_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_J_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_K_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // JKFFSRXL
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFSX1 (Q, QN, VDD, VSS, CK, J, K, SN);
inout VDD, VSS;
output Q, QN;
input  J, K, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;
  buf   XX0 (xSN, SN);

udp_jkff_PWR  I0 (n0,J, K,CK,xRN,xSN,VDD, VSS, NOTIFIER); 
buf I1 (Q,n0);
not I2 (QN,n0);

wire ENABLE_J_AND_SN_OR_K_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_K ;
assign ENABLE_J_AND_SN_OR_K_AND_SN = (J&SN | K&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_K = (K) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_J_AND_SN_OR_K_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_J_AND_SN_OR_K_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_K == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // JKFFSX1
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFSX2 (Q, QN, VDD, VSS, CK, J, K, SN);
inout VDD, VSS;
output Q, QN;
input  J, K, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;
  buf   XX0 (xSN, SN);

udp_jkff_PWR  I0 (n0,J, K,CK,xRN,xSN,VDD, VSS, NOTIFIER); 
buf I1 (Q,n0);
not I2 (QN,n0);

wire ENABLE_J_AND_SN_OR_K_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_K ;
assign ENABLE_J_AND_SN_OR_K_AND_SN = (J&SN | K&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_K = (K) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_J_AND_SN_OR_K_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_J_AND_SN_OR_K_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_K == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // JKFFSX2
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFSX4 (Q, QN, VDD, VSS, CK, J, K, SN);
inout VDD, VSS;
output Q, QN;
input  J, K, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;
  buf   XX0 (xSN, SN);

udp_jkff_PWR  I0 (n0,J, K,CK,xRN,xSN,VDD, VSS, NOTIFIER); 
buf I1 (Q,n0);
not I2 (QN,n0);

wire ENABLE_J_AND_SN_OR_K_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_K ;
assign ENABLE_J_AND_SN_OR_K_AND_SN = (J&SN | K&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_K = (K) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_J_AND_SN_OR_K_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_J_AND_SN_OR_K_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_K == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // JKFFSX4
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFSXL (Q, QN, VDD, VSS, CK, J, K, SN);
inout VDD, VSS;
output Q, QN;
input  J, K, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;
  buf   XX0 (xSN, SN);

udp_jkff_PWR  I0 (n0,J, K,CK,xRN,xSN,VDD, VSS, NOTIFIER); 
buf I1 (Q,n0);
not I2 (QN,n0);

wire ENABLE_J_AND_SN_OR_K_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_K ;
assign ENABLE_J_AND_SN_OR_K_AND_SN = (J&SN | K&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_K = (K) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_J_AND_SN_OR_K_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_J_AND_SN_OR_K_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_K == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // JKFFSXL
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFX1 (Q, QN, VDD, VSS, CK, J, K);
inout VDD, VSS;
output Q, QN;
input  J, K, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

udp_jkff_PWR  I0 (n0,J, K,CK,xRN,xSN,VDD, VSS, NOTIFIER); 
buf I1 (Q,n0);
not I2 (QN,n0);

wire ENABLE_J_OR_K ;
assign ENABLE_J_OR_K = (J | K) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_J_OR_K == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_J_OR_K == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, posedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // JKFFX1
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFX2 (Q, QN, VDD, VSS, CK, J, K);
inout VDD, VSS;
output Q, QN;
input  J, K, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

udp_jkff_PWR  I0 (n0,J, K,CK,xRN,xSN,VDD, VSS, NOTIFIER); 
buf I1 (Q,n0);
not I2 (QN,n0);

wire ENABLE_J_OR_K ;
assign ENABLE_J_OR_K = (J | K) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_J_OR_K == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_J_OR_K == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, posedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // JKFFX2
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFX4 (Q, QN, VDD, VSS, CK, J, K);
inout VDD, VSS;
output Q, QN;
input  J, K, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

udp_jkff_PWR  I0 (n0,J, K,CK,xRN,xSN,VDD, VSS, NOTIFIER); 
buf I1 (Q,n0);
not I2 (QN,n0);

wire ENABLE_J_OR_K ;
assign ENABLE_J_OR_K = (J | K) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_J_OR_K == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_J_OR_K == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, posedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // JKFFX4
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFXL (Q, QN, VDD, VSS, CK, J, K);
inout VDD, VSS;
output Q, QN;
input  J, K, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

udp_jkff_PWR  I0 (n0,J, K,CK,xRN,xSN,VDD, VSS, NOTIFIER); 
buf I1 (Q,n0);
not I2 (QN,n0);

wire ENABLE_J_OR_K ;
assign ENABLE_J_OR_K = (J | K) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_J_OR_K == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_J_OR_K == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, posedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // JKFFXL
`endcelldefine





`timescale 1ns/1ps
`celldefine
module MX2X1 (Y, VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2X2 (Y, VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2X4 (Y, VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2XL (Y, VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(out_temp, A, B, S0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX4X1 (Y, VDD, VSS, A, B, C, D, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(out_temp, A, B, C, D, S0, S1);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX4X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX4X2 (Y, VDD, VSS, A, B, C, D, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(out_temp, A, B, C, D, S0, S1);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX4X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX4X4 (Y, VDD, VSS, A, B, C, D, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(out_temp, A, B, C, D, S0, S1);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX4X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX4XL (Y, VDD, VSS, A, B, C, D, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(out_temp, A, B, C, D, S0, S1);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX4XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2X1 (Y, VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI2X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2X2 (Y, VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI2X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2X4 (Y, VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI2X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2XL (Y, VDD, VSS, A, B, S0);
inout VDD, VSS;
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI2XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI4X1 (Y, VDD, VSS, A, B, C, D, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI4X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI4X2 (Y, VDD, VSS, A, B, C, D, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI4X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI4X4 (Y, VDD, VSS, A, B, C, D, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI4X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI4XL (Y, VDD, VSS, A, B, C, D, S0, S1);
inout VDD, VSS;
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(out_temp, YN);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI4XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2BX1 (Y, VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nand (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2BX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2BX2 (Y, VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nand (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2BX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2BX4 (Y, VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nand (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2BX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2BXL (Y, VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nand (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2BXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2X1 (Y, VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2X2 (Y, VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2X4 (Y, VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2XL (Y, VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nand (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BX1 (Y, VDD, VSS, AN, B, C);
inout VDD, VSS;
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (out_temp, Ax, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3BX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BX2 (Y, VDD, VSS, AN, B, C);
inout VDD, VSS;
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (out_temp, Ax, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3BX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BX4 (Y, VDD, VSS, AN, B, C);
inout VDD, VSS;
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (out_temp, Ax, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3BX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BXL (Y, VDD, VSS, AN, B, C);
inout VDD, VSS;
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (out_temp, Ax, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3BXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3X1 (Y, VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nand (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3X2 (Y, VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nand (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3X4 (Y, VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nand (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3XL (Y, VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nand (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BBX1 (Y, VDD, VSS, AN, BN, C, D);
inout VDD, VSS;
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (out_temp, Ax, Bx, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BBX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BBX2 (Y, VDD, VSS, AN, BN, C, D);
inout VDD, VSS;
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (out_temp, Ax, Bx, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BBX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BBX4 (Y, VDD, VSS, AN, BN, C, D);
inout VDD, VSS;
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (out_temp, Ax, Bx, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BBX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BBXL (Y, VDD, VSS, AN, BN, C, D);
inout VDD, VSS;
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (out_temp, Ax, Bx, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BBXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BX1 (Y, VDD, VSS, AN, B, C, D);
inout VDD, VSS;
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (out_temp, Ax, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BX2 (Y, VDD, VSS, AN, B, C, D);
inout VDD, VSS;
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (out_temp, Ax, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BX4 (Y, VDD, VSS, AN, B, C, D);
inout VDD, VSS;
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (out_temp, Ax, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BXL (Y, VDD, VSS, AN, B, C, D);
inout VDD, VSS;
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (out_temp, Ax, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4X1 (Y, VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nand (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4X2 (Y, VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nand (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4X4 (Y, VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nand (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4XL (Y, VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nand (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2BX1 (Y, VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nor (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2BX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2BX2 (Y, VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nor (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2BX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2BX4 (Y, VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nor (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2BX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2BXL (Y, VDD, VSS, AN, B);
inout VDD, VSS;
output Y;
input AN, B;

  not (Ax, AN);
  nor (out_temp, Ax, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2BXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2X1 (Y, VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2X2 (Y, VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2X4 (Y, VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2XL (Y, VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  nor (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BX1 (Y, VDD, VSS, AN, B, C);
inout VDD, VSS;
output Y;
input AN, B, C;

  not (Ax, AN);
  nor (out_temp, Ax, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3BX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BX2 (Y, VDD, VSS, AN, B, C);
inout VDD, VSS;
output Y;
input AN, B, C;

  not (Ax, AN);
  nor (out_temp, Ax, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3BX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BX4 (Y, VDD, VSS, AN, B, C);
inout VDD, VSS;
output Y;
input AN, B, C;

  not (Ax, AN);
  nor (out_temp, Ax, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3BX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BXL (Y, VDD, VSS, AN, B, C);
inout VDD, VSS;
output Y;
input AN, B, C;

  not (Ax, AN);
  nor (out_temp, Ax, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3BXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3X1 (Y, VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nor (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3X2 (Y, VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nor (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3X4 (Y, VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nor (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3XL (Y, VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  nor (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BBX1 (Y, VDD, VSS, AN, BN, C, D);
inout VDD, VSS;
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor (out_temp, Ax, Bx, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BBX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BBX2 (Y, VDD, VSS, AN, BN, C, D);
inout VDD, VSS;
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor (out_temp, Ax, Bx, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BBX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BBX4 (Y, VDD, VSS, AN, BN, C, D);
inout VDD, VSS;
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor (out_temp, Ax, Bx, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BBX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BBXL (Y, VDD, VSS, AN, BN, C, D);
inout VDD, VSS;
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor (out_temp, Ax, Bx, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BBXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BX1 (Y, VDD, VSS, AN, B, C, D);
inout VDD, VSS;
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nor (out_temp, Ax, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BX2 (Y, VDD, VSS, AN, B, C, D);
inout VDD, VSS;
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nor (out_temp, Ax, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BX4 (Y, VDD, VSS, AN, B, C, D);
inout VDD, VSS;
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nor (out_temp, Ax, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BXL (Y, VDD, VSS, AN, B, C, D);
inout VDD, VSS;
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nor (out_temp, Ax, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4X1 (Y, VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nor (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4X2 (Y, VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nor (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4X4 (Y, VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nor (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4XL (Y, VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  nor (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211X1 (Y, VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI211X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211X2 (Y, VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI211X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211X4 (Y, VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI211X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211XL (Y, VDD, VSS, A0, A1, B0, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, C0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI211XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21X1 (Y, VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21X2 (Y, VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21X4 (Y, VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21XL (Y, VDD, VSS, A0, A1, B0);
inout VDD, VSS;
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221X1 (Y, VDD, VSS, A0, A1, B0, B1, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(out_temp, C0, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI221X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221X2 (Y, VDD, VSS, A0, A1, B0, B1, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(out_temp, C0, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI221X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221X4 (Y, VDD, VSS, A0, A1, B0, B1, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(out_temp, C0, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI221X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221XL (Y, VDD, VSS, A0, A1, B0, B1, C0);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(out_temp, C0, outB, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI221XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222X1 (Y, VDD, VSS, A0, A1, B0, B1, C0, C1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(out_temp, outA, outB, outC);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI222X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222X2 (Y, VDD, VSS, A0, A1, B0, B1, C0, C1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(out_temp, outA, outB, outC);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI222X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222X4 (Y, VDD, VSS, A0, A1, B0, B1, C0, C1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(out_temp, outA, outB, outC);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI222X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222XL (Y, VDD, VSS, A0, A1, B0, B1, C0, C1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(out_temp, outA, outB, outC);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI222XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22X1 (Y, VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22X2 (Y, VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22X4 (Y, VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22XL (Y, VDD, VSS, A0, A1, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB1X1 (Y, VDD, VSS, A0N, A1N, B0);
inout VDD, VSS;
output Y;
input A0N, A1N, B0;



  nand I0 (outA, A0N, A1N);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2BB1X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB1X2 (Y, VDD, VSS, A0N, A1N, B0);
inout VDD, VSS;
output Y;
input A0N, A1N, B0;



  nand I0 (outA, A0N, A1N);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2BB1X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB1X4 (Y, VDD, VSS, A0N, A1N, B0);
inout VDD, VSS;
output Y;
input A0N, A1N, B0;



  nand I0 (outA, A0N, A1N);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2BB1X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB1XL (Y, VDD, VSS, A0N, A1N, B0);
inout VDD, VSS;
output Y;
input A0N, A1N, B0;



  nand I0 (outA, A0N, A1N);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2BB1XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB2X1 (Y, VDD, VSS, A0N, A1N, B0, B1);
inout VDD, VSS;
output Y;
input A0N, A1N, B0, B1;



  nand I0 (outA, A0N, A1N);
  or   I1(outB, B0, B1);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2BB2X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB2X2 (Y, VDD, VSS, A0N, A1N, B0, B1);
inout VDD, VSS;
output Y;
input A0N, A1N, B0, B1;



  nand I0 (outA, A0N, A1N);
  or   I1(outB, B0, B1);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2BB2X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB2X4 (Y, VDD, VSS, A0N, A1N, B0, B1);
inout VDD, VSS;
output Y;
input A0N, A1N, B0, B1;



  nand I0 (outA, A0N, A1N);
  or   I1(outB, B0, B1);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2BB2X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB2XL (Y, VDD, VSS, A0N, A1N, B0, B1);
inout VDD, VSS;
output Y;
input A0N, A1N, B0, B1;



  nand I0 (outA, A0N, A1N);
  or   I1(outB, B0, B1);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2BB2XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31X1 (Y, VDD, VSS, A0, A1, A2, B0);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI31X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31X2 (Y, VDD, VSS, A0, A1, A2, B0);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI31X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31X4 (Y, VDD, VSS, A0, A1, A2, B0);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI31X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31XL (Y, VDD, VSS, A0, A1, A2, B0);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand I1(out_temp, B0, outA);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI31XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI32X1 (Y, VDD, VSS, A0, A1, A2, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI32X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI32X2 (Y, VDD, VSS, A0, A1, A2, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI32X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI32X4 (Y, VDD, VSS, A0, A1, A2, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI32X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI32XL (Y, VDD, VSS, A0, A1, A2, B0, B1);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI32XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI33X1 (Y, VDD, VSS, A0, A1, A2, B0, B1, B2);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1, B2;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1, B2);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI33X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI33X2 (Y, VDD, VSS, A0, A1, A2, B0, B1, B2);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1, B2;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1, B2);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI33X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI33X4 (Y, VDD, VSS, A0, A1, A2, B0, B1, B2);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1, B2;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1, B2);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI33X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI33XL (Y, VDD, VSS, A0, A1, A2, B0, B1, B2);
inout VDD, VSS;
output Y;
input A0, A1, A2, B0, B1, B2;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1, B2);
  nand I2(out_temp, outA, outB);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI33XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2X1 (Y, VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  or (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2X2 (Y, VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  or (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2X4 (Y, VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  or (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2XL (Y, VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  or (out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3X1 (Y, VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  or (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3X2 (Y, VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  or (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3X4 (Y, VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  or (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3XL (Y, VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  or (out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4X1 (Y, VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  or (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4X2 (Y, VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  or (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4X4 (Y, VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  or (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4XL (Y, VDD, VSS, A, B, C, D);
inout VDD, VSS;
output Y;
input A, B, C, D;

  or (out_temp, A, B, C, D);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF1R1WX2 (RB, VDD, VSS, RW, RWN, WB, WW);
inout VDD, VSS;
output RB;
input WB, WW, RW, RWN;
reg NOTIFIER;

   not II (wwn,WW);
   udp_tlatrf_PWR  I0 (n0, WB, WW, wwn, VDD, VSS, NOTIFIER);
   notif1     I1 (rdbl_temp, n0, n2);
  assign RB = ((VDD === 1'b1) && (VSS === 1'b0))? rdbl_temp : 1'bx;
   udp_outrf  I2 (n2, n0, RWN, RW);





wire ENABLE_RW_AND_NOT_RWN ;
assign ENABLE_RW_AND_NOT_RWN = (RW&!RWN) ? 1'b1:1'b0;

specify
(WB => RB) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WB==1'b0 && WW==1'b0)
( RW => RB ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WB==1'b1 && WW==1'b0)
( RW => RB ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WW==1'b1)
( RW => RB ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WB==1'b0 && WW==1'b0)
( RWN => RB ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WB==1'b1 && WW==1'b0)
( RWN => RB ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WW==1'b1)
( RWN => RB ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge WW &&& (ENABLE_RW_AND_NOT_RWN == 1'b1), posedge WB, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WW &&& (ENABLE_RW_AND_NOT_RWN == 1'b1), negedge WB, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge WW &&& (ENABLE_RW_AND_NOT_RWN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge WW => (RB:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // RF1R1WX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF2R1WX2 (R1B, R2B, VDD, VSS, R1W, R2W, WB, WW);
inout VDD, VSS;
output R1B, R2B;
input WB, WW, R1W, R2W;
reg NOTIFIER;

   not        I0 (WWN, WW);
   not        I1 (R1WN, R1W);
   not        I2 (R2WN, R2W);
   udp_tlatrf_PWR  I3 (n0, WB, WW, WWN, VDD, VSS, NOTIFIER);
   notif1     I4 (rdbl1_temp, n0, n2);
  assign R1B = ((VDD === 1'b1) && (VSS === 1'b0))? rdbl1_temp : 1'bx;
   notif1     I5 (rdbl2_temp, n0, n3);
  assign R2B = ((VDD === 1'b1) && (VSS === 1'b0))? rdbl2_temp : 1'bx;
   udp_outrf  I6 (n2, n0, R1WN, R1W);
   udp_outrf  I7 (n3, n0, R2WN, R2W);





wire ENABLE_R1W_OR_R2W ;
assign ENABLE_R1W_OR_R2W = (R1W | R2W) ? 1'b1:1'b0;

specify
if (R2W==1'b0)
(WB => R1B) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R2W==1'b1)
(WB => R1B) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R1W==1'b0)
(WB => R2B) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R1W==1'b1)
(WB => R2B) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R2W==1'b0 && WB==1'b0 && WW==1'b0)
( R1W => R1B ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R2W==1'b0 && WB==1'b1 && WW==1'b0)
( R1W => R1B ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R2W==1'b0 && WW==1'b1)
( R1W => R1B ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R2W==1'b1 && WB==1'b0 && WW==1'b0)
( R1W => R1B ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R2W==1'b1 && WB==1'b1 && WW==1'b0)
( R1W => R1B ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R2W==1'b1 && WW==1'b1)
( R1W => R1B ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R1W==1'b0 && WB==1'b0 && WW==1'b0)
( R2W => R2B ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R1W==1'b0 && WB==1'b1 && WW==1'b0)
( R2W => R2B ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R1W==1'b0 && WW==1'b1)
( R2W => R2B ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R1W==1'b1 && WB==1'b0 && WW==1'b0)
( R2W => R2B ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R1W==1'b1 && WB==1'b1 && WW==1'b0)
( R2W => R2B ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R1W==1'b1 && WW==1'b1)
( R2W => R2B ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge WW &&& (ENABLE_R1W_OR_R2W == 1'b1), posedge WB, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WW &&& (ENABLE_R1W_OR_R2W == 1'b1), negedge WB, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge WW &&& (ENABLE_R1W_OR_R2W == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (R2W==1'b0)
(posedge WW => (R1B:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R2W==1'b1)
(posedge WW => (R1B:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R1W==1'b0)
(posedge WW => (R2B:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R1W==1'b1)
(posedge WW => (R2B:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // RF2R1WX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RFRDX1 (BRB, VDD, VSS, RB);
inout VDD, VSS;
output BRB;
input RB;
reg NOTIFIER;

   not(weak0,weak1) I0(RB, io_wire);
   not              I1(io_wire, RB);
   buf              I2(out_temp, io_wire);
  assign BRB = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;






specify
(RB => BRB) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // RFRDX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RFRDX2 (BRB, VDD, VSS, RB);
inout VDD, VSS;
output BRB;
input RB;
reg NOTIFIER;

   not(weak0,weak1) I0(RB, io_wire);
   not              I1(io_wire, RB);
   buf              I2(out_temp, io_wire);
  assign BRB = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;






specify
(RB => BRB) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // RFRDX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RFRDX4 (BRB, VDD, VSS, RB);
inout VDD, VSS;
output BRB;
input RB;
reg NOTIFIER;

   not(weak0,weak1) I0(RB, io_wire);
   not              I1(io_wire, RB);
   buf              I2(out_temp, io_wire);
  assign BRB = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;






specify
(RB => BRB) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // RFRDX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RSLATNX1 (Q, QN, VDD, VSS, RN, SN);
inout VDD, VSS;
output Q, QN;
input RN, SN;
reg NOTIFIER;
  not I4(R, RN);
  not I5(S, SN);
  udp_rslat_pwr  I0(q,  R, S, VDD, VSS, NOTIFIER);
  udp_rslatn_pwr I1(qn, R, S, VDD, VSS, NOTIFIER);
  not I2(QN, q);
  not I3(Q, qn);

wire ENABLE_SN ;
wire ENABLE_RN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge SN, posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (SN==1'b0)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (SN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // RSLATNX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RSLATNX2 (Q, QN, VDD, VSS, RN, SN);
inout VDD, VSS;
output Q, QN;
input RN, SN;
reg NOTIFIER;
  not I4(R, RN);
  not I5(S, SN);
  udp_rslat_pwr  I0(q,  R, S, VDD, VSS, NOTIFIER);
  udp_rslatn_pwr I1(qn, R, S, VDD, VSS, NOTIFIER);
  not I2(QN, q);
  not I3(Q, qn);

wire ENABLE_SN ;
wire ENABLE_RN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge SN, posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (SN==1'b0)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (SN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // RSLATNX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RSLATNX4 (Q, QN, VDD, VSS, RN, SN);
inout VDD, VSS;
output Q, QN;
input RN, SN;
reg NOTIFIER;
  not I4(R, RN);
  not I5(S, SN);
  udp_rslat_pwr  I0(q,  R, S, VDD, VSS, NOTIFIER);
  udp_rslatn_pwr I1(qn, R, S, VDD, VSS, NOTIFIER);
  not I2(QN, q);
  not I3(Q, qn);

wire ENABLE_SN ;
wire ENABLE_RN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge SN, posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (SN==1'b0)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (SN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // RSLATNX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RSLATNXL (Q, QN, VDD, VSS, RN, SN);
inout VDD, VSS;
output Q, QN;
input RN, SN;
reg NOTIFIER;
  not I4(R, RN);
  not I5(S, SN);
  udp_rslat_pwr  I0(q,  R, S, VDD, VSS, NOTIFIER);
  udp_rslatn_pwr I1(qn, R, S, VDD, VSS, NOTIFIER);
  not I2(QN, q);
  not I3(Q, qn);

wire ENABLE_SN ;
wire ENABLE_RN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge SN, posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (SN==1'b0)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (SN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // RSLATNXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RSLATX1 (Q, QN, VDD, VSS, R, S);
inout VDD, VSS;
output Q, QN;
input R, S;
reg NOTIFIER;
  udp_rslat_pwr  I0(q, R, S, VDD, VSS, NOTIFIER);
  udp_rslatn_pwr  I1(qn, R, S, VDD, VSS, NOTIFIER);
  buf I2(QN, qn);
  buf I3(Q, q);


wire ENABLE_NOT_S ;
wire ENABLE_NOT_R ;
assign ENABLE_NOT_S = (!S) ? 1'b1:1'b0;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;

specify
$width(posedge R &&& (ENABLE_NOT_S == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge S, negedge R, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R, negedge S, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge S &&& (ENABLE_NOT_R == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (S==1'b0)
(posedge R *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (S==1'b1)
(R => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (R==1'b0)
(posedge S *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (R==1'b1)
(S => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // RSLATX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RSLATX2 (Q, QN, VDD, VSS, R, S);
inout VDD, VSS;
output Q, QN;
input R, S;
reg NOTIFIER;
  udp_rslat_pwr  I0(q, R, S, VDD, VSS, NOTIFIER);
  udp_rslatn_pwr  I1(qn, R, S, VDD, VSS, NOTIFIER);
  buf I2(QN, qn);
  buf I3(Q, q);


wire ENABLE_NOT_S ;
wire ENABLE_NOT_R ;
assign ENABLE_NOT_S = (!S) ? 1'b1:1'b0;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;

specify
$width(posedge R &&& (ENABLE_NOT_S == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge S, negedge R, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R, negedge S, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge S &&& (ENABLE_NOT_R == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (S==1'b0)
(posedge R *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (S==1'b1)
(R => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (R==1'b0)
(posedge S *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (R==1'b1)
(S => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // RSLATX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RSLATX4 (Q, QN, VDD, VSS, R, S);
inout VDD, VSS;
output Q, QN;
input R, S;
reg NOTIFIER;
  udp_rslat_pwr  I0(q, R, S, VDD, VSS, NOTIFIER);
  udp_rslatn_pwr  I1(qn, R, S, VDD, VSS, NOTIFIER);
  buf I2(QN, qn);
  buf I3(Q, q);


wire ENABLE_NOT_S ;
wire ENABLE_NOT_R ;
assign ENABLE_NOT_S = (!S) ? 1'b1:1'b0;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;

specify
$width(posedge R &&& (ENABLE_NOT_S == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge S, negedge R, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R, negedge S, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge S &&& (ENABLE_NOT_R == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (S==1'b0)
(posedge R *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (S==1'b1)
(R => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (R==1'b0)
(posedge S *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (R==1'b1)
(S => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // RSLATX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RSLATXL (Q, QN, VDD, VSS, R, S);
inout VDD, VSS;
output Q, QN;
input R, S;
reg NOTIFIER;
  udp_rslat_pwr  I0(q, R, S, VDD, VSS, NOTIFIER);
  udp_rslatn_pwr  I1(qn, R, S, VDD, VSS, NOTIFIER);
  buf I2(QN, qn);
  buf I3(Q, q);


wire ENABLE_NOT_S ;
wire ENABLE_NOT_R ;
assign ENABLE_NOT_S = (!S) ? 1'b1:1'b0;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;

specify
$width(posedge R &&& (ENABLE_NOT_S == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge S, negedge R, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R, negedge S, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge S &&& (ENABLE_NOT_R == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (S==1'b0)
(posedge R *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (S==1'b1)
(R => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (R==1'b0)
(posedge S *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (R==1'b1)
(S => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // RSLATXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module SDFFHQX1 (Q, VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI = (D&!SI | !D&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFHQX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFHQX2 (Q, VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI = (D&!SI | !D&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFHQX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFHQX4 (Q, VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI = (D&!SI | !D&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFHQX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFHQXL (Q, VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI = (D&!SI | !D&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFHQXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNRX1 (Q, QN, VDD, VSS, CKN, D, RN, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CKN, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  not     IC (clk, CKN);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI = (D&!SE | SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI = (D&RN&!SI | !D&RN&SI) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, negedge CKN &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // SDFFNRX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNRX2 (Q, QN, VDD, VSS, CKN, D, RN, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CKN, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  not     IC (clk, CKN);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI = (D&!SE | SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI = (D&RN&!SI | !D&RN&SI) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, negedge CKN &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // SDFFNRX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNRX4 (Q, QN, VDD, VSS, CKN, D, RN, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CKN, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  not     IC (clk, CKN);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI = (D&!SE | SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI = (D&RN&!SI | !D&RN&SI) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, negedge CKN &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // SDFFNRX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNRXL (Q, QN, VDD, VSS, CKN, D, RN, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CKN, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  not     IC (clk, CKN);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI = (D&!SE | SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI = (D&RN&!SI | !D&RN&SI) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, negedge CKN &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // SDFFNRXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSRX1 (Q, QN, VDD, VSS, CKN, D, RN, SE, SI, SN);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CKN, SN, RN;
reg NOTIFIER;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN = (D&!SE&SN | SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN = (D&RN&!SI&SN | !D&RN&SI&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI = (!D&RN&!SE | RN&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNSRX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSRX2 (Q, QN, VDD, VSS, CKN, D, RN, SE, SI, SN);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CKN, SN, RN;
reg NOTIFIER;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN = (D&!SE&SN | SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN = (D&RN&!SI&SN | !D&RN&SI&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI = (!D&RN&!SE | RN&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNSRX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSRX4 (Q, QN, VDD, VSS, CKN, D, RN, SE, SI, SN);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CKN, SN, RN;
reg NOTIFIER;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN = (D&!SE&SN | SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN = (D&RN&!SI&SN | !D&RN&SI&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI = (!D&RN&!SE | RN&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNSRX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSRXL (Q, QN, VDD, VSS, CKN, D, RN, SE, SI, SN);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CKN, SN, RN;
reg NOTIFIER;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN = (D&!SE&SN | SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN = (D&RN&!SI&SN | !D&RN&SI&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI = (!D&RN&!SE | RN&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNSRXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSX1 (Q, QN, VDD, VSS, CKN, D, SE, SI, SN);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CKN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN ;
wire ENABLE_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN = (D&!SI&SN | !D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI = (!D&!SE | SE&!SI) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNSX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSX2 (Q, QN, VDD, VSS, CKN, D, SE, SI, SN);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CKN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN ;
wire ENABLE_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN = (D&!SI&SN | !D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI = (!D&!SE | SE&!SI) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNSX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSX4 (Q, QN, VDD, VSS, CKN, D, SE, SI, SN);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CKN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN ;
wire ENABLE_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN = (D&!SI&SN | !D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI = (!D&!SE | SE&!SI) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNSX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSXL (Q, QN, VDD, VSS, CKN, D, SE, SI, SN);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CKN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN ;
wire ENABLE_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN = (D&!SI&SN | !D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI = (!D&!SE | SE&!SI) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNSXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNX1 (Q, QN, VDD, VSS, CKN, D, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CKN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, CKN);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI = (D&!SI | !D&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CKN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFNX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNX2 (Q, QN, VDD, VSS, CKN, D, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CKN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, CKN);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI = (D&!SI | !D&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CKN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFNX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNX4 (Q, QN, VDD, VSS, CKN, D, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CKN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, CKN);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI = (D&!SI | !D&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CKN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFNX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNXL (Q, QN, VDD, VSS, CKN, D, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CKN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, CKN);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI = (D&!SI | !D&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CKN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFNXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRHQX1 (Q, VDD, VSS, CK, D, RN, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI = (D&!SE | SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI = (D&RN&!SI | !D&RN&SI) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFRHQX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRHQX2 (Q, VDD, VSS, CK, D, RN, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI = (D&!SE | SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI = (D&RN&!SI | !D&RN&SI) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFRHQX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRHQX4 (Q, VDD, VSS, CK, D, RN, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI = (D&!SE | SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI = (D&RN&!SI | !D&RN&SI) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFRHQX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRHQXL (Q, VDD, VSS, CK, D, RN, SE, SI);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI = (D&!SE | SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI = (D&RN&!SI | !D&RN&SI) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFRHQXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRX1 (Q, QN, VDD, VSS, CK, D, RN, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI = (D&!SE | SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI = (D&RN&!SI | !D&RN&SI) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // SDFFRX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRX2 (Q, QN, VDD, VSS, CK, D, RN, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI = (D&!SE | SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI = (D&RN&!SI | !D&RN&SI) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // SDFFRX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRX4 (Q, QN, VDD, VSS, CK, D, RN, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI = (D&!SE | SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI = (D&RN&!SI | !D&RN&SI) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // SDFFRX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRXL (Q, QN, VDD, VSS, CK, D, RN, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI = (D&!SE | SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI = (D&RN&!SI | !D&RN&SI) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // SDFFRXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSHQX1 (Q, VDD, VSS, CK, D, SE, SI, SN);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN ;
wire ENABLE_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN = (D&!SI&SN | !D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI = (!D&!SE | SE&!SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // SDFFSHQX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSHQX2 (Q, VDD, VSS, CK, D, SE, SI, SN);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN ;
wire ENABLE_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN = (D&!SI&SN | !D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI = (!D&!SE | SE&!SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // SDFFSHQX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSHQX4 (Q, VDD, VSS, CK, D, SE, SI, SN);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN ;
wire ENABLE_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN = (D&!SI&SN | !D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI = (!D&!SE | SE&!SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // SDFFSHQX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSHQXL (Q, VDD, VSS, CK, D, SE, SI, SN);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN ;
wire ENABLE_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN = (D&!SI&SN | !D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI = (!D&!SE | SE&!SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // SDFFSHQXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRHQX1 (Q, VDD, VSS, CK, D, RN, SE, SI, SN);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN = (D&!SE&SN | SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN = (D&RN&!SI&SN | !D&RN&SI&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI = (!D&RN&!SE | RN&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // SDFFSRHQX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRHQX2 (Q, VDD, VSS, CK, D, RN, SE, SI, SN);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN = (D&!SE&SN | SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN = (D&RN&!SI&SN | !D&RN&SI&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI = (!D&RN&!SE | RN&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // SDFFSRHQX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRHQX4 (Q, VDD, VSS, CK, D, RN, SE, SI, SN);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN = (D&!SE&SN | SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN = (D&RN&!SI&SN | !D&RN&SI&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI = (!D&RN&!SE | RN&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // SDFFSRHQX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRHQXL (Q, VDD, VSS, CK, D, RN, SE, SI, SN);
inout VDD, VSS;
output Q;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN = (D&!SE&SN | SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN = (D&RN&!SI&SN | !D&RN&SI&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI = (!D&RN&!SE | RN&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // SDFFSRHQXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRX1 (Q, QN, VDD, VSS, CK, D, RN, SE, SI, SN);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN = (D&!SE&SN | SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN = (D&RN&!SI&SN | !D&RN&SI&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI = (!D&RN&!SE | RN&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSRX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRX2 (Q, QN, VDD, VSS, CK, D, RN, SE, SI, SN);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN = (D&!SE&SN | SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN = (D&RN&!SI&SN | !D&RN&SI&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI = (!D&RN&!SE | RN&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSRX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRX4 (Q, QN, VDD, VSS, CK, D, RN, SE, SI, SN);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN = (D&!SE&SN | SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN = (D&RN&!SI&SN | !D&RN&SI&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI = (!D&RN&!SE | RN&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSRX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRXL (Q, QN, VDD, VSS, CK, D, RN, SE, SI, SN);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN = (D&!SE&SN | SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN = (D&RN&!SI&SN | !D&RN&SI&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI = (!D&RN&!SE | RN&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSRXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSX1 (Q, QN, VDD, VSS, CK, D, SE, SI, SN);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN ;
wire ENABLE_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN = (D&!SI&SN | !D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI = (!D&!SE | SE&!SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSX2 (Q, QN, VDD, VSS, CK, D, SE, SI, SN);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN ;
wire ENABLE_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN = (D&!SI&SN | !D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI = (!D&!SE | SE&!SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSX4 (Q, QN, VDD, VSS, CK, D, SE, SI, SN);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN ;
wire ENABLE_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN = (D&!SI&SN | !D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI = (!D&!SE | SE&!SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSXL (Q, QN, VDD, VSS, CK, D, SE, SI, SN);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN ;
wire ENABLE_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN = (D&!SI&SN | !D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI = (!D&!SE | SE&!SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFTRX1 (Q, QN, VDD, VSS, CK, D, RN, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
   udp_sedfft_PWR  I0 (n0, D, CK, xRN, SI, SE, 1'b1, VDD, VSS, NOTIFIER);
   buf        I1 (Q, n0);
   not        I2 (QN, n0);

wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_RN_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE = (D&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_RN_AND_SI = (D&RN&!SI | !D&SI | !RN&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFTRX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFTRX2 (Q, QN, VDD, VSS, CK, D, RN, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
   udp_sedfft_PWR  I0 (n0, D, CK, xRN, SI, SE, 1'b1, VDD, VSS, NOTIFIER);
   buf        I1 (Q, n0);
   not        I2 (QN, n0);

wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_RN_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE = (D&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_RN_AND_SI = (D&RN&!SI | !D&SI | !RN&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFTRX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFTRX4 (Q, QN, VDD, VSS, CK, D, RN, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
   udp_sedfft_PWR  I0 (n0, D, CK, xRN, SI, SE, 1'b1, VDD, VSS, NOTIFIER);
   buf        I1 (Q, n0);
   not        I2 (QN, n0);

wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_RN_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE = (D&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_RN_AND_SI = (D&RN&!SI | !D&SI | !RN&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFTRX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFTRXL (Q, QN, VDD, VSS, CK, D, RN, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
   udp_sedfft_PWR  I0 (n0, D, CK, xRN, SI, SE, 1'b1, VDD, VSS, NOTIFIER);
   buf        I1 (Q, n0);
   not        I2 (QN, n0);

wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_RN_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE = (D&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_RN_AND_SI = (D&RN&!SI | !D&SI | !RN&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFTRXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFX1 (Q, QN, VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI = (D&!SI | !D&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFX2 (Q, QN, VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI = (D&!SI | !D&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFX4 (Q, QN, VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI = (D&!SI | !D&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFXL (Q, QN, VDD, VSS, CK, D, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff_PWR  I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI = (D&!SI | !D&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SEDFFHQX1 (Q, VDD, VSS, CK, D, E, SE, SI);
inout VDD, VSS;
output Q;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR  I0 (n0, D, CK, xRN, SI, SE, E, VDD, VSS, NOTIFIER);
   buf       I1 (Q, n0);

wire ENABLE_E_OR_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E ;
wire ENABLE_SE ;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E = (D&!SI | !D&SI | !E) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFHQX1
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFHQX2 (Q, VDD, VSS, CK, D, E, SE, SI);
inout VDD, VSS;
output Q;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR  I0 (n0, D, CK, xRN, SI, SE, E, VDD, VSS, NOTIFIER);
   buf       I1 (Q, n0);

wire ENABLE_E_OR_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E ;
wire ENABLE_SE ;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E = (D&!SI | !D&SI | !E) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFHQX2
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFHQX4 (Q, VDD, VSS, CK, D, E, SE, SI);
inout VDD, VSS;
output Q;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR  I0 (n0, D, CK, xRN, SI, SE, E, VDD, VSS, NOTIFIER);
   buf       I1 (Q, n0);

wire ENABLE_E_OR_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E ;
wire ENABLE_SE ;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E = (D&!SI | !D&SI | !E) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFHQX4
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFHQXL (Q, VDD, VSS, CK, D, E, SE, SI);
inout VDD, VSS;
output Q;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR  I0 (n0, D, CK, xRN, SI, SE, E, VDD, VSS, NOTIFIER);
   buf       I1 (Q, n0);

wire ENABLE_E_OR_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E ;
wire ENABLE_SE ;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E = (D&!SI | !D&SI | !E) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFHQXL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFTRX1 (Q, QN, VDD, VSS, CK, D, E, RN, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, CK, E, SE, SI, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

   udp_sedfft_PWR  I0 (n0, D, CK, xRN, SI, SE, E, VDD, VSS, NOTIFIER);
   buf        I1 (Q, n0);
   not        I2 (QN, n0);

wire ENABLE_E_OR_NOT_RN_OR_SE ;
wire ENABLE_E_AND_RN_AND_NOT_SE ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE_OR_NOT_E_AND_NOT_SE ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E_AND_RN_OR_NOT_RN_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_E_OR_NOT_RN_OR_SE = (E | !RN | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_RN_AND_NOT_SE = (E&RN&!SE) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_OR_NOT_E_AND_NOT_SE = (D&!SE | !E&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E_AND_RN_OR_NOT_RN_AND_SI = (D&RN&!SI | !D&SI | !E&RN | !RN&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_NOT_RN_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_NOT_RN_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_NOT_E_AND_NOT_SE == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_NOT_E_AND_NOT_SE == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E_AND_RN_OR_NOT_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E_AND_RN_OR_NOT_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFTRX1
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFTRX2 (Q, QN, VDD, VSS, CK, D, E, RN, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, CK, E, SE, SI, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

   udp_sedfft_PWR  I0 (n0, D, CK, xRN, SI, SE, E, VDD, VSS, NOTIFIER);
   buf        I1 (Q, n0);
   not        I2 (QN, n0);

wire ENABLE_E_OR_NOT_RN_OR_SE ;
wire ENABLE_E_AND_RN_AND_NOT_SE ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE_OR_NOT_E_AND_NOT_SE ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E_AND_RN_OR_NOT_RN_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_E_OR_NOT_RN_OR_SE = (E | !RN | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_RN_AND_NOT_SE = (E&RN&!SE) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_OR_NOT_E_AND_NOT_SE = (D&!SE | !E&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E_AND_RN_OR_NOT_RN_AND_SI = (D&RN&!SI | !D&SI | !E&RN | !RN&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_NOT_RN_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_NOT_RN_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_NOT_E_AND_NOT_SE == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_NOT_E_AND_NOT_SE == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E_AND_RN_OR_NOT_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E_AND_RN_OR_NOT_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFTRX2
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFTRX4 (Q, QN, VDD, VSS, CK, D, E, RN, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, CK, E, SE, SI, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

   udp_sedfft_PWR  I0 (n0, D, CK, xRN, SI, SE, E, VDD, VSS, NOTIFIER);
   buf        I1 (Q, n0);
   not        I2 (QN, n0);

wire ENABLE_E_OR_NOT_RN_OR_SE ;
wire ENABLE_E_AND_RN_AND_NOT_SE ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE_OR_NOT_E_AND_NOT_SE ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E_AND_RN_OR_NOT_RN_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_E_OR_NOT_RN_OR_SE = (E | !RN | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_RN_AND_NOT_SE = (E&RN&!SE) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_OR_NOT_E_AND_NOT_SE = (D&!SE | !E&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E_AND_RN_OR_NOT_RN_AND_SI = (D&RN&!SI | !D&SI | !E&RN | !RN&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_NOT_RN_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_NOT_RN_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_NOT_E_AND_NOT_SE == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_NOT_E_AND_NOT_SE == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E_AND_RN_OR_NOT_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E_AND_RN_OR_NOT_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFTRX4
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFTRXL (Q, QN, VDD, VSS, CK, D, E, RN, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, CK, E, SE, SI, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

   udp_sedfft_PWR  I0 (n0, D, CK, xRN, SI, SE, E, VDD, VSS, NOTIFIER);
   buf        I1 (Q, n0);
   not        I2 (QN, n0);

wire ENABLE_E_OR_NOT_RN_OR_SE ;
wire ENABLE_E_AND_RN_AND_NOT_SE ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE_OR_NOT_E_AND_NOT_SE ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E_AND_RN_OR_NOT_RN_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_E_OR_NOT_RN_OR_SE = (E | !RN | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_RN_AND_NOT_SE = (E&RN&!SE) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_OR_NOT_E_AND_NOT_SE = (D&!SE | !E&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E_AND_RN_OR_NOT_RN_AND_SI = (D&RN&!SI | !D&SI | !E&RN | !RN&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_NOT_RN_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_NOT_RN_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_NOT_E_AND_NOT_SE == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_NOT_E_AND_NOT_SE == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E_AND_RN_OR_NOT_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E_AND_RN_OR_NOT_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFTRXL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFX1 (Q, QN, VDD, VSS, CK, D, E, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR  I0 (n0, D, CK, xRN, SI, SE, E, VDD, VSS, NOTIFIER); 
  buf     I1 (Q, n0);  
  not     I2 (QN, n0);

wire ENABLE_E_OR_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E ;
wire ENABLE_SE ;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E = (D&!SI | !D&SI | !E) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFX1
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFX2 (Q, QN, VDD, VSS, CK, D, E, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR  I0 (n0, D, CK, xRN, SI, SE, E, VDD, VSS, NOTIFIER); 
  buf     I1 (Q, n0);  
  not     I2 (QN, n0);

wire ENABLE_E_OR_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E ;
wire ENABLE_SE ;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E = (D&!SI | !D&SI | !E) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFX2
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFX4 (Q, QN, VDD, VSS, CK, D, E, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR  I0 (n0, D, CK, xRN, SI, SE, E, VDD, VSS, NOTIFIER); 
  buf     I1 (Q, n0);  
  not     I2 (QN, n0);

wire ENABLE_E_OR_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E ;
wire ENABLE_SE ;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E = (D&!SI | !D&SI | !E) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFX4
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFXL (Q, QN, VDD, VSS, CK, D, E, SE, SI);
inout VDD, VSS;
output Q, QN;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR  I0 (n0, D, CK, xRN, SI, SE, E, VDD, VSS, NOTIFIER); 
  buf     I1 (Q, n0);  
  not     I2 (QN, n0);

wire ENABLE_E_OR_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E ;
wire ENABLE_SE ;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E = (D&!SI | !D&SI | !E) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFXL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module TBUFIX1 (Y, VDD, VSS, A, OE);
inout VDD, VSS;
output Y;
input A, OE;

  notif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFIX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFIX12 (Y, VDD, VSS, A, OE);
inout VDD, VSS;
output Y;
input A, OE;

  notif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFIX12
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFIX16 (Y, VDD, VSS, A, OE);
inout VDD, VSS;
output Y;
input A, OE;

  notif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFIX16
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFIX2 (Y, VDD, VSS, A, OE);
inout VDD, VSS;
output Y;
input A, OE;

  notif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFIX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFIX20 (Y, VDD, VSS, A, OE);
inout VDD, VSS;
output Y;
input A, OE;

  notif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFIX20
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFIX3 (Y, VDD, VSS, A, OE);
inout VDD, VSS;
output Y;
input A, OE;

  notif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFIX3
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFIX4 (Y, VDD, VSS, A, OE);
inout VDD, VSS;
output Y;
input A, OE;

  notif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFIX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFIX8 (Y, VDD, VSS, A, OE);
inout VDD, VSS;
output Y;
input A, OE;

  notif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFIX8
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFIXL (Y, VDD, VSS, A, OE);
inout VDD, VSS;
output Y;
input A, OE;

  notif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFIXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFX1 (Y, VDD, VSS, A, OE);
inout VDD, VSS;
output Y;
input A, OE;

  bufif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFX12 (Y, VDD, VSS, A, OE);
inout VDD, VSS;
output Y;
input A, OE;

  bufif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFX12
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFX16 (Y, VDD, VSS, A, OE);
inout VDD, VSS;
output Y;
input A, OE;

  bufif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFX16
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFX2 (Y, VDD, VSS, A, OE);
inout VDD, VSS;
output Y;
input A, OE;

  bufif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFX20 (Y, VDD, VSS, A, OE);
inout VDD, VSS;
output Y;
input A, OE;

  bufif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFX20
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFX3 (Y, VDD, VSS, A, OE);
inout VDD, VSS;
output Y;
input A, OE;

  bufif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFX3
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFX4 (Y, VDD, VSS, A, OE);
inout VDD, VSS;
output Y;
input A, OE;

  bufif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFX8 (Y, VDD, VSS, A, OE);
inout VDD, VSS;
output Y;
input A, OE;

  bufif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFX8
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFXL (Y, VDD, VSS, A, OE);
inout VDD, VSS;
output Y;
input A, OE;

  bufif1 I0(out_temp, A, OE);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TIEHI (Y, VDD, VSS);
inout VDD, VSS;
output Y;

  buf I0(out_temp, 1'b1);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify

endspecify
endmodule // TIEHI
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TIELO (Y, VDD, VSS);
inout VDD, VSS;
output Y;

  buf I0(out_temp, 1'b0);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


specify

endspecify
endmodule // TIELO
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATCOX1 (ECKN, VDD, VSS, CKN, E);
inout VDD, VSS;
output ECKN;
input  E, CKN;
reg NOTIFIER;

supply1 R, S;

  not      I0 (nclk,CKN);
  udp_tlat_PWR  I1 (n0, E, nclk, R, S, VDD, VSS, NOTIFIER);
  not      I2 (nn0,n0);
  or       I3 (out_temp, nn0, CKN);
  assign ECKN = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CKN => ECKN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(posedge CKN => (ECKN:1'bx)) = (`ARM_PROP_DELAY,`ARM_INVALID_DELAY);
$width(posedge CKN &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(posedge CKN &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATCOX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATCOX2 (ECKN, VDD, VSS, CKN, E);
inout VDD, VSS;
output ECKN;
input  E, CKN;
reg NOTIFIER;

supply1 R, S;

  not      I0 (nclk,CKN);
  udp_tlat_PWR  I1 (n0, E, nclk, R, S, VDD, VSS, NOTIFIER);
  not      I2 (nn0,n0);
  or       I3 (out_temp, nn0, CKN);
  assign ECKN = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CKN => ECKN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(posedge CKN => (ECKN:1'bx)) = (`ARM_PROP_DELAY,`ARM_INVALID_DELAY);
$width(posedge CKN &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(posedge CKN &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATCOX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATCOX3 (ECKN, VDD, VSS, CKN, E);
inout VDD, VSS;
output ECKN;
input  E, CKN;
reg NOTIFIER;

supply1 R, S;

  not      I0 (nclk,CKN);
  udp_tlat_PWR  I1 (n0, E, nclk, R, S, VDD, VSS, NOTIFIER);
  not      I2 (nn0,n0);
  or       I3 (out_temp, nn0, CKN);
  assign ECKN = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CKN => ECKN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(posedge CKN => (ECKN:1'bx)) = (`ARM_PROP_DELAY,`ARM_INVALID_DELAY);
$width(posedge CKN &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(posedge CKN &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATCOX3
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATCOX4 (ECKN, VDD, VSS, CKN, E);
inout VDD, VSS;
output ECKN;
input  E, CKN;
reg NOTIFIER;

supply1 R, S;

  not      I0 (nclk,CKN);
  udp_tlat_PWR  I1 (n0, E, nclk, R, S, VDD, VSS, NOTIFIER);
  not      I2 (nn0,n0);
  or       I3 (out_temp, nn0, CKN);
  assign ECKN = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CKN => ECKN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(posedge CKN => (ECKN:1'bx)) = (`ARM_PROP_DELAY,`ARM_INVALID_DELAY);
$width(posedge CKN &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(posedge CKN &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATCOX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNCAX1 (ECK, VDD, VSS, CK, E);
inout VDD, VSS;
output ECK;
input  E, CK;
reg NOTIFIER;

supply1 R, S;

  udp_tlat_PWR  I0 (n0, E, CK, R, S, VDD, VSS, NOTIFIER);
  and      I1 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(negedge CK => (ECK:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATNCAX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNCAX2 (ECK, VDD, VSS, CK, E);
inout VDD, VSS;
output ECK;
input  E, CK;
reg NOTIFIER;

supply1 R, S;

  udp_tlat_PWR  I0 (n0, E, CK, R, S, VDD, VSS, NOTIFIER);
  and      I1 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(negedge CK => (ECK:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATNCAX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNCAX3 (ECK, VDD, VSS, CK, E);
inout VDD, VSS;
output ECK;
input  E, CK;
reg NOTIFIER;

supply1 R, S;

  udp_tlat_PWR  I0 (n0, E, CK, R, S, VDD, VSS, NOTIFIER);
  and      I1 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(negedge CK => (ECK:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATNCAX3
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNCAX4 (ECK, VDD, VSS, CK, E);
inout VDD, VSS;
output ECK;
input  E, CK;
reg NOTIFIER;

supply1 R, S;

  udp_tlat_PWR  I0 (n0, E, CK, R, S, VDD, VSS, NOTIFIER);
  and      I1 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(negedge CK => (ECK:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATNCAX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNCAX6 (ECK, VDD, VSS, CK, E);
inout VDD, VSS;
output ECK;
input  E, CK;
reg NOTIFIER;

supply1 R, S;

  udp_tlat_PWR  I0 (n0, E, CK, R, S, VDD, VSS, NOTIFIER);
  and      I1 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(negedge CK => (ECK:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATNCAX6
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNCAX8 (ECK, VDD, VSS, CK, E);
inout VDD, VSS;
output ECK;
input  E, CK;
reg NOTIFIER;

supply1 R, S;

  udp_tlat_PWR  I0 (n0, E, CK, R, S, VDD, VSS, NOTIFIER);
  and      I1 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(negedge CK => (ECK:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATNCAX8
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNRX1 (Q, QN, VDD, VSS, D, GN, RN);
inout VDD, VSS;
output  Q, QN;
input  D, GN, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);
udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, GN);

wire ENABLE_RN ;
wire ENABLE_D ;
wire ENABLE_GN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_GN = (GN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge RN, posedge GN &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_GN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // TLATNRX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNRX2 (Q, QN, VDD, VSS, D, GN, RN);
inout VDD, VSS;
output  Q, QN;
input  D, GN, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);
udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, GN);

wire ENABLE_RN ;
wire ENABLE_D ;
wire ENABLE_GN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_GN = (GN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge RN, posedge GN &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_GN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // TLATNRX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNRX4 (Q, QN, VDD, VSS, D, GN, RN);
inout VDD, VSS;
output  Q, QN;
input  D, GN, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);
udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, GN);

wire ENABLE_RN ;
wire ENABLE_D ;
wire ENABLE_GN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_GN = (GN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge RN, posedge GN &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_GN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // TLATNRX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNRXL (Q, QN, VDD, VSS, D, GN, RN);
inout VDD, VSS;
output  Q, QN;
input  D, GN, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);
udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, GN);

wire ENABLE_RN ;
wire ENABLE_D ;
wire ENABLE_GN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_GN = (GN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge RN, posedge GN &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_GN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // TLATNRXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNSRX1 (Q, QN, VDD, VSS, D, GN, RN, SN);
inout VDD, VSS;
output  Q, QN;
input  D, GN, RN, SN;
reg NOTIFIER;

buf       XX0 (xSN, SN);
buf       XX1 (xRN, RN);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_GN_AND_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_GN ;
wire ENABLE_GN_AND_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_GN_AND_SN = (GN&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_GN = (GN) ? 1'b1:1'b0;
assign ENABLE_GN_AND_RN = (GN&RN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge RN, posedge GN &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_GN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge GN &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN &&& (ENABLE_GN == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_GN_AND_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && GN==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATNSRX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNSRX2 (Q, QN, VDD, VSS, D, GN, RN, SN);
inout VDD, VSS;
output  Q, QN;
input  D, GN, RN, SN;
reg NOTIFIER;

buf       XX0 (xSN, SN);
buf       XX1 (xRN, RN);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_GN_AND_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_GN ;
wire ENABLE_GN_AND_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_GN_AND_SN = (GN&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_GN = (GN) ? 1'b1:1'b0;
assign ENABLE_GN_AND_RN = (GN&RN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge RN, posedge GN &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_GN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge GN &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN &&& (ENABLE_GN == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_GN_AND_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && GN==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATNSRX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNSRX4 (Q, QN, VDD, VSS, D, GN, RN, SN);
inout VDD, VSS;
output  Q, QN;
input  D, GN, RN, SN;
reg NOTIFIER;

buf       XX0 (xSN, SN);
buf       XX1 (xRN, RN);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_GN_AND_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_GN ;
wire ENABLE_GN_AND_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_GN_AND_SN = (GN&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_GN = (GN) ? 1'b1:1'b0;
assign ENABLE_GN_AND_RN = (GN&RN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge RN, posedge GN &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_GN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge GN &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN &&& (ENABLE_GN == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_GN_AND_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && GN==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATNSRX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNSRXL (Q, QN, VDD, VSS, D, GN, RN, SN);
inout VDD, VSS;
output  Q, QN;
input  D, GN, RN, SN;
reg NOTIFIER;

buf       XX0 (xSN, SN);
buf       XX1 (xRN, RN);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_GN_AND_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_GN ;
wire ENABLE_GN_AND_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_GN_AND_SN = (GN&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_GN = (GN) ? 1'b1:1'b0;
assign ENABLE_GN_AND_RN = (GN&RN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge RN, posedge GN &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_GN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge GN &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN &&& (ENABLE_GN == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_GN_AND_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && GN==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATNSRXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNSX1 (Q, QN, VDD, VSS, D, GN, SN);
inout VDD, VSS;
output  Q, QN;
input  D, GN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);
udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, GN);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_GN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_GN = (GN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_GN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATNSX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNSX2 (Q, QN, VDD, VSS, D, GN, SN);
inout VDD, VSS;
output  Q, QN;
input  D, GN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);
udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, GN);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_GN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_GN = (GN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_GN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATNSX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNSX4 (Q, QN, VDD, VSS, D, GN, SN);
inout VDD, VSS;
output  Q, QN;
input  D, GN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);
udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, GN);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_GN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_GN = (GN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_GN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATNSX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNSXL (Q, QN, VDD, VSS, D, GN, SN);
inout VDD, VSS;
output  Q, QN;
input  D, GN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);
udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, GN);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_GN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_GN = (GN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_GN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATNSXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNTSCAX1 (ECK, VDD, VSS, CK, E, SE);
inout VDD, VSS;
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR  I1 (n0, n1, CK, R, S, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATNTSCAX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNTSCAX2 (ECK, VDD, VSS, CK, E, SE);
inout VDD, VSS;
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR  I1 (n0, n1, CK, R, S, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATNTSCAX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNTSCAX3 (ECK, VDD, VSS, CK, E, SE);
inout VDD, VSS;
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR  I1 (n0, n1, CK, R, S, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATNTSCAX3
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNTSCAX4 (ECK, VDD, VSS, CK, E, SE);
inout VDD, VSS;
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR  I1 (n0, n1, CK, R, S, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATNTSCAX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNTSCAX6 (ECK, VDD, VSS, CK, E, SE);
inout VDD, VSS;
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR  I1 (n0, n1, CK, R, S, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATNTSCAX6
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNTSCAX8 (ECK, VDD, VSS, CK, E, SE);
inout VDD, VSS;
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR  I1 (n0, n1, CK, R, S, VDD, VSS, NOTIFIER);
  and      I2 (out_temp, n0, CK);
  assign ECK = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATNTSCAX8
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNX1 (Q, QN, VDD, VSS, D, GN);
inout VDD, VSS;
output  Q, QN;
input  D, GN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);


specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TLATNX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNX2 (Q, QN, VDD, VSS, D, GN);
inout VDD, VSS;
output  Q, QN;
input  D, GN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);


specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TLATNX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNX4 (Q, QN, VDD, VSS, D, GN);
inout VDD, VSS;
output  Q, QN;
input  D, GN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);


specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TLATNX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNXL (Q, QN, VDD, VSS, D, GN);
inout VDD, VSS;
output  Q, QN;
input  D, GN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);


specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TLATNXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATRX1 (Q, QN, VDD, VSS, D, G, RN);
inout VDD, VSS;
output  Q, QN;
input  D, G, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);
udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_RN ;
wire ENABLE_D ;
wire ENABLE_NOT_G ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_G = (!G) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge RN, negedge G &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_NOT_G == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b1)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATRX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATRX2 (Q, QN, VDD, VSS, D, G, RN);
inout VDD, VSS;
output  Q, QN;
input  D, G, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);
udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_RN ;
wire ENABLE_D ;
wire ENABLE_NOT_G ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_G = (!G) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge RN, negedge G &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_NOT_G == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b1)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATRX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATRX4 (Q, QN, VDD, VSS, D, G, RN);
inout VDD, VSS;
output  Q, QN;
input  D, G, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);
udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_RN ;
wire ENABLE_D ;
wire ENABLE_NOT_G ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_G = (!G) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge RN, negedge G &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_NOT_G == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b1)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATRX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATRXL (Q, QN, VDD, VSS, D, G, RN);
inout VDD, VSS;
output  Q, QN;
input  D, G, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);
udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_RN ;
wire ENABLE_D ;
wire ENABLE_NOT_G ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_G = (!G) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge RN, negedge G &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_NOT_G == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b1)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATRXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATSRX1 (Q, QN, VDD, VSS, D, G, RN, SN);
inout VDD, VSS;
output  Q, QN;
input  D, G, SN, RN;
reg NOTIFIER;

buf       XX0 (xSN, SN);
buf       XX1 (xRN, RN);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_G_AND_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_NOT_G ;
wire ENABLE_NOT_G_AND_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_G_AND_SN = (!G&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_NOT_G = (!G) ? 1'b1:1'b0;
assign ENABLE_NOT_G_AND_RN = (!G&RN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge RN, negedge G &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_NOT_G_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, negedge G &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN &&& (ENABLE_NOT_G == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_G_AND_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b1)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATSRX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATSRX2 (Q, QN, VDD, VSS, D, G, RN, SN);
inout VDD, VSS;
output  Q, QN;
input  D, G, SN, RN;
reg NOTIFIER;

buf       XX0 (xSN, SN);
buf       XX1 (xRN, RN);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_G_AND_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_NOT_G ;
wire ENABLE_NOT_G_AND_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_G_AND_SN = (!G&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_NOT_G = (!G) ? 1'b1:1'b0;
assign ENABLE_NOT_G_AND_RN = (!G&RN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge RN, negedge G &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_NOT_G_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, negedge G &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN &&& (ENABLE_NOT_G == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_G_AND_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b1)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATSRX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATSRX4 (Q, QN, VDD, VSS, D, G, RN, SN);
inout VDD, VSS;
output  Q, QN;
input  D, G, SN, RN;
reg NOTIFIER;

buf       XX0 (xSN, SN);
buf       XX1 (xRN, RN);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_G_AND_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_NOT_G ;
wire ENABLE_NOT_G_AND_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_G_AND_SN = (!G&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_NOT_G = (!G) ? 1'b1:1'b0;
assign ENABLE_NOT_G_AND_RN = (!G&RN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge RN, negedge G &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_NOT_G_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, negedge G &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN &&& (ENABLE_NOT_G == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_G_AND_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b1)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATSRX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATSRXL (Q, QN, VDD, VSS, D, G, RN, SN);
inout VDD, VSS;
output  Q, QN;
input  D, G, SN, RN;
reg NOTIFIER;

buf       XX0 (xSN, SN);
buf       XX1 (xRN, RN);

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_G_AND_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_NOT_G ;
wire ENABLE_NOT_G_AND_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_G_AND_SN = (!G&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_NOT_G = (!G) ? 1'b1:1'b0;
assign ENABLE_NOT_G_AND_RN = (!G&RN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge RN, negedge G &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_NOT_G_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, negedge G &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN &&& (ENABLE_NOT_G == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_G_AND_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b1)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATSRXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATSX1 (Q, QN, VDD, VSS, D, G, SN);
inout VDD, VSS;
output  Q, QN;
input  D, G, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);
udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_G ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_G = (!G) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, negedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_G == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && G==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATSX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATSX2 (Q, QN, VDD, VSS, D, G, SN);
inout VDD, VSS;
output  Q, QN;
input  D, G, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);
udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_G ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_G = (!G) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, negedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_G == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && G==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATSX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATSX4 (Q, QN, VDD, VSS, D, G, SN);
inout VDD, VSS;
output  Q, QN;
input  D, G, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);
udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_G ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_G = (!G) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, negedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_G == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && G==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATSX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATSXL (Q, QN, VDD, VSS, D, G, SN);
inout VDD, VSS;
output  Q, QN;
input  D, G, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);
udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_G ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_G = (!G) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, negedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_G == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && G==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATSXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATTSCOX1 (ECKN, VDD, VSS, CKN, E, SE);
inout VDD, VSS;
output ECKN;
input  E, SE, CKN;
reg NOTIFIER;

supply1 R, S;

  not      I0 (nclk,CKN);
  or       I1 (n1, SE, E);
  udp_tlat_PWR  I2 (n0, n1, nclk, R, S, VDD, VSS, NOTIFIER);
  not      I3 (nn0,n0);
  or       I4 (out_temp, nn0, CKN);
  assign ECKN = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CKN => ECKN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CKN => ECKN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CKN => ECKN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(posedge CKN => (ECKN:1'bx)) = (`ARM_PROP_DELAY,`ARM_INVALID_DELAY);
$width(posedge CKN &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(posedge CKN &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATTSCOX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATTSCOX2 (ECKN, VDD, VSS, CKN, E, SE);
inout VDD, VSS;
output ECKN;
input  E, SE, CKN;
reg NOTIFIER;

supply1 R, S;

  not      I0 (nclk,CKN);
  or       I1 (n1, SE, E);
  udp_tlat_PWR  I2 (n0, n1, nclk, R, S, VDD, VSS, NOTIFIER);
  not      I3 (nn0,n0);
  or       I4 (out_temp, nn0, CKN);
  assign ECKN = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CKN => ECKN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CKN => ECKN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CKN => ECKN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(posedge CKN => (ECKN:1'bx)) = (`ARM_PROP_DELAY,`ARM_INVALID_DELAY);
$width(posedge CKN &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(posedge CKN &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATTSCOX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATTSCOX3 (ECKN, VDD, VSS, CKN, E, SE);
inout VDD, VSS;
output ECKN;
input  E, SE, CKN;
reg NOTIFIER;

supply1 R, S;

  not      I0 (nclk,CKN);
  or       I1 (n1, SE, E);
  udp_tlat_PWR  I2 (n0, n1, nclk, R, S, VDD, VSS, NOTIFIER);
  not      I3 (nn0,n0);
  or       I4 (out_temp, nn0, CKN);
  assign ECKN = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CKN => ECKN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CKN => ECKN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CKN => ECKN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(posedge CKN => (ECKN:1'bx)) = (`ARM_PROP_DELAY,`ARM_INVALID_DELAY);
$width(posedge CKN &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(posedge CKN &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATTSCOX3
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATTSCOX4 (ECKN, VDD, VSS, CKN, E, SE);
inout VDD, VSS;
output ECKN;
input  E, SE, CKN;
reg NOTIFIER;

supply1 R, S;

  not      I0 (nclk,CKN);
  or       I1 (n1, SE, E);
  udp_tlat_PWR  I2 (n0, n1, nclk, R, S, VDD, VSS, NOTIFIER);
  not      I3 (nn0,n0);
  or       I4 (out_temp, nn0, CKN);
  assign ECKN = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CKN => ECKN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CKN => ECKN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CKN => ECKN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(posedge CKN => (ECKN:1'bx)) = (`ARM_PROP_DELAY,`ARM_INVALID_DELAY);
$width(posedge CKN &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(posedge CKN &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATTSCOX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATX1 (Q, QN, VDD, VSS, D, G);
inout VDD, VSS;
output  Q, QN;
input  D, G;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,G);


specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TLATX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATX2 (Q, QN, VDD, VSS, D, G);
inout VDD, VSS;
output  Q, QN;
input  D, G;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,G);


specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TLATX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATX4 (Q, QN, VDD, VSS, D, G);
inout VDD, VSS;
output  Q, QN;
input  D, G;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,G);


specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TLATX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATXL (Q, QN, VDD, VSS, D, G);
inout VDD, VSS;
output  Q, QN;
input  D, G;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,G);


specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TLATXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TTLATX1 (Q, VDD, VSS, D, G, OE);
inout VDD, VSS;
output Q;
input  D, G, OE;
reg NOTIFIER;
supply1 RN, SN;
supply1 xRN, xSN;
supply1 dRN, dSN;

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
bufif1   I1 (out_temp, n0, OE);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
not  I3(clk,G);

wire ENABLE_OE ;
assign ENABLE_OE = (OE) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
( OE => Q ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
( OE => Q ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (G==1'b1)
( OE => Q ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_OE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_OE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_OE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TTLATX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TTLATX2 (Q, VDD, VSS, D, G, OE);
inout VDD, VSS;
output Q;
input  D, G, OE;
reg NOTIFIER;
supply1 RN, SN;
supply1 xRN, xSN;
supply1 dRN, dSN;

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
bufif1   I1 (out_temp, n0, OE);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
not  I3(clk,G);

wire ENABLE_OE ;
assign ENABLE_OE = (OE) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
( OE => Q ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
( OE => Q ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (G==1'b1)
( OE => Q ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_OE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_OE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_OE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TTLATX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TTLATX4 (Q, VDD, VSS, D, G, OE);
inout VDD, VSS;
output Q;
input  D, G, OE;
reg NOTIFIER;
supply1 RN, SN;
supply1 xRN, xSN;
supply1 dRN, dSN;

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
bufif1   I1 (out_temp, n0, OE);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
not  I3(clk,G);

wire ENABLE_OE ;
assign ENABLE_OE = (OE) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
( OE => Q ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
( OE => Q ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (G==1'b1)
( OE => Q ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_OE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_OE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_OE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TTLATX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TTLATXL (Q, VDD, VSS, D, G, OE);
inout VDD, VSS;
output Q;
input  D, G, OE;
reg NOTIFIER;
supply1 RN, SN;
supply1 xRN, xSN;
supply1 dRN, dSN;

udp_tlat_PWR  I0 (n0, D, clk, xRN, xSN, VDD, VSS, NOTIFIER);
bufif1   I1 (out_temp, n0, OE);
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;
not  I3(clk,G);

wire ENABLE_OE ;
assign ENABLE_OE = (OE) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
( OE => Q ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
( OE => Q ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (G==1'b1)
( OE => Q ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_OE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_OE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_OE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TTLATXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2X1 (Y, VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xnor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR2X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2X2 (Y, VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xnor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR2X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2X4 (Y, VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xnor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR2X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2XL (Y, VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xnor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR2XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3X2 (Y, VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  xnor I0(out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR3X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3X4 (Y, VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  xnor I0(out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR3X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2X1 (Y, VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR2X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2X2 (Y, VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR2X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2X4 (Y, VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR2X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2XL (Y, VDD, VSS, A, B);
inout VDD, VSS;
output Y;
input A, B;

  xor I0(out_temp, A, B);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR2XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3X2 (Y, VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  xor I0(out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR3X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3X4 (Y, VDD, VSS, A, B, C);
inout VDD, VSS;
output Y;
input A, B, C;

  xor I0(out_temp, A, B, C);
  assign Y = ((VDD === 1'b1) && (VSS === 1'b0))? out_temp : 1'bx;



specify
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR3X4
`endcelldefine
`else

`timescale 1ns/1ps
`celldefine
module ADDFHX1 (CO, S, A, B, CI);
output S, CO;
input A, B, CI;
  xor I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFHX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFHX2 (CO, S, A, B, CI);
output S, CO;
input A, B, CI;
  xor I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFHX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFHX4 (CO, S, A, B, CI);
output S, CO;
input A, B, CI;
  xor I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFHX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFHXL (CO, S, A, B, CI);
output S, CO;
input A, B, CI;
  xor I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFHXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFX1 (CO, S, A, B, CI);
output S, CO;
input A, B, CI;
  xor I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFX2 (CO, S, A, B, CI);
output S, CO;
input A, B, CI;
  xor I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFX4 (CO, S, A, B, CI);
output S, CO;
input A, B, CI;
  xor I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDFXL (CO, S, A, B, CI);
output S, CO;
input A, B, CI;
  xor I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or I4(CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDFXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDHX1 (CO, S, A, B);
output S, CO;
input A, B;
  xor I0(S, A, B);
  and I1(CO, A, B);


specify
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDHX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDHX2 (CO, S, A, B);
output S, CO;
input A, B;
  xor I0(S, A, B);
  and I1(CO, A, B);


specify
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDHX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDHX4 (CO, S, A, B);
output S, CO;
input A, B;
  xor I0(S, A, B);
  and I1(CO, A, B);


specify
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDHX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ADDHXL (CO, S, A, B);
output S, CO;
input A, B;
  xor I0(S, A, B);
  and I1(CO, A, B);


specify
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // ADDHXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AFCSHCINX2 (CO0, CO1, S, A, B, CI0N, CI1N, CS);
output S, CO0, CO1;
input A, B, CI0N, CI1N, CS;
  not I0 (cin1, CI1N);
  not I1 (cin0, CI0N);
  xor I2 (s1, A, B, cin1);
  xor I3 (s2, A, B, cin0);
  and I4 (s3, CS, s1);
  not I5 (csn, CS);
  and I6 (s4, csn, s2);
  or I7 (S, s3, s4);
  and I8 (a_and_b, A, B);
  and I9 (a_and_ci0, A, cin0);
  and I10 (b_and_ci0, B, cin0);
  or I11 (CO0, a_and_b, a_and_ci0, b_and_ci0);
  and I12 (a_and_ci1, A, cin1);
  and I13 (b_and_ci1, B, cin1);
  or I14 (CO1, a_and_b, a_and_ci1, b_and_ci1);


specify
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b0)
(A => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b1)
(A => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b0)
(A => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b1)
(A => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b0)
(A => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b1)
(A => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b0)
(A => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b1)
(A => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b0)
(B => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b1)
(B => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b0)
(B => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b1)
(B => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b0)
(B => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b1)
(B => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b0)
(B => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b1)
(B => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1N==1'b0 && CS==1'b0)
(CI0N => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1N==1'b0 && CS==1'b1)
(CI0N => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1N==1'b1 && CS==1'b0)
(CI0N => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1N==1'b1 && CS==1'b1)
(CI0N => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1N==1'b0 && CS==1'b0)
(CI0N => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1N==1'b0 && CS==1'b1)
(CI0N => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1N==1'b1 && CS==1'b0)
(CI0N => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1N==1'b1 && CS==1'b1)
(CI0N => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b0)
(A => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b1)
(A => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b0)
(A => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b1)
(A => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b0)
(A => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b1)
(A => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b0)
(A => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b1)
(A => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b0)
(B => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b1)
(B => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b0)
(B => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b1)
(B => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b0)
(B => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b1)
(B => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b0)
(B => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b1)
(B => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0N==1'b0 && CS==1'b0)
(CI1N => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0N==1'b0 && CS==1'b1)
(CI1N => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0N==1'b1 && CS==1'b0)
(CI1N => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0N==1'b1 && CS==1'b1)
(CI1N => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0N==1'b0 && CS==1'b0)
(CI1N => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0N==1'b0 && CS==1'b1)
(CI1N => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0N==1'b1 && CS==1'b0)
(CI1N => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0N==1'b1 && CS==1'b1)
(CI1N => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI1N==1'b0)
(CI0N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI1N==1'b1)
(CI0N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI1N==1'b0)
(CI0N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI1N==1'b1)
(CI0N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1N==1'b0)
(CI0N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1N==1'b1)
(CI0N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1N==1'b0)
(CI0N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1N==1'b1)
(CI0N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI0N==1'b0)
(CI1N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI0N==1'b1)
(CI1N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI0N==1'b0)
(CI1N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI0N==1'b1)
(CI1N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0N==1'b0)
(CI1N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0N==1'b1)
(CI1N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0N==1'b0)
(CI1N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0N==1'b1)
(CI1N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI0N==1'b0 && CI1N==1'b1)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0N==1'b1 && CI1N==1'b0)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0N==1'b1 && CI1N==1'b0)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI0N==1'b0 && CI1N==1'b1)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI0N==1'b1 && CI1N==1'b0)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0N==1'b0 && CI1N==1'b1)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0N==1'b0 && CI1N==1'b1)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI0N==1'b1 && CI1N==1'b0)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AFCSHCINX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AFCSHCINX4 (CO0, CO1, S, A, B, CI0N, CI1N, CS);
output S, CO0, CO1;
input A, B, CI0N, CI1N, CS;
  not I0 (cin1, CI1N);
  not I1 (cin0, CI0N);
  xor I2 (s1, A, B, cin1);
  xor I3 (s2, A, B, cin0);
  and I4 (s3, CS, s1);
  not I5 (csn, CS);
  and I6 (s4, csn, s2);
  or I7 (S, s3, s4);
  and I8 (a_and_b, A, B);
  and I9 (a_and_ci0, A, cin0);
  and I10 (b_and_ci0, B, cin0);
  or I11 (CO0, a_and_b, a_and_ci0, b_and_ci0);
  and I12 (a_and_ci1, A, cin1);
  and I13 (b_and_ci1, B, cin1);
  or I14 (CO1, a_and_b, a_and_ci1, b_and_ci1);


specify
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b0)
(A => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b1)
(A => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b0)
(A => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b1)
(A => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b0)
(A => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b1)
(A => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b0)
(A => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b1)
(A => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b0)
(B => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b1)
(B => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b0)
(B => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b1)
(B => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b0)
(B => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b1)
(B => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b0)
(B => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b1)
(B => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1N==1'b0 && CS==1'b0)
(CI0N => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1N==1'b0 && CS==1'b1)
(CI0N => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1N==1'b1 && CS==1'b0)
(CI0N => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1N==1'b1 && CS==1'b1)
(CI0N => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1N==1'b0 && CS==1'b0)
(CI0N => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1N==1'b0 && CS==1'b1)
(CI0N => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1N==1'b1 && CS==1'b0)
(CI0N => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1N==1'b1 && CS==1'b1)
(CI0N => CO0) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b0)
(A => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b1)
(A => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b0)
(A => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b1)
(A => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b0)
(A => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b1)
(A => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b0)
(A => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b1)
(A => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b0)
(B => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b1)
(B => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b0)
(B => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b1)
(B => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b0)
(B => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b1)
(B => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b0)
(B => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b1)
(B => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0N==1'b0 && CS==1'b0)
(CI1N => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0N==1'b0 && CS==1'b1)
(CI1N => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0N==1'b1 && CS==1'b0)
(CI1N => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0N==1'b1 && CS==1'b1)
(CI1N => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0N==1'b0 && CS==1'b0)
(CI1N => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0N==1'b0 && CS==1'b1)
(CI1N => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0N==1'b1 && CS==1'b0)
(CI1N => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0N==1'b1 && CS==1'b1)
(CI1N => CO1) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0N==1'b1 && CI1N==1'b1 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b0 && CI1N==1'b0 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b0 && CI1N==1'b1 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0N==1'b1 && CI1N==1'b0 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI1N==1'b0)
(CI0N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI1N==1'b1)
(CI0N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI1N==1'b0)
(CI0N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI1N==1'b1)
(CI0N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1N==1'b0)
(CI0N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1N==1'b1)
(CI0N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1N==1'b0)
(CI0N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1N==1'b1)
(CI0N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI0N==1'b0)
(CI1N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI0N==1'b1)
(CI1N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI0N==1'b0)
(CI1N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI0N==1'b1)
(CI1N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0N==1'b0)
(CI1N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0N==1'b1)
(CI1N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0N==1'b0)
(CI1N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0N==1'b1)
(CI1N => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI0N==1'b0 && CI1N==1'b1)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0N==1'b1 && CI1N==1'b0)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0N==1'b1 && CI1N==1'b0)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI0N==1'b0 && CI1N==1'b1)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI0N==1'b1 && CI1N==1'b0)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0N==1'b0 && CI1N==1'b1)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0N==1'b0 && CI1N==1'b1)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI0N==1'b1 && CI1N==1'b0)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AFCSHCINX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AFCSHCONX2 (CO0N, CO1N, S, A, B, CI0, CI1, CS);
output S, CO0N, CO1N;
input A, B, CI0, CI1, CS;
  xor I2 (s1, A, B, CI1);
  xor I3 (s2, A, B, CI0);
  and I4 (s3, CS, s1);
  not I5 (csn, CS);
  and I6 (s4, csn, s2);
  or I7 (S, s3, s4);
  and I8 (a_and_b, A, B);
  and I9 (a_and_ci0, A, CI0);
  and I10 (b_and_ci0, B, CI0);
  or I11 (cout0, a_and_b, a_and_ci0, b_and_ci0);
  and I12 (a_and_ci1, A, CI1);
  and I13 (b_and_ci1, B, CI1);
  or I14 (cout1, a_and_b, a_and_ci1, b_and_ci1);
  not I15 (CO0N, cout0);
  not I16 (CO1N, cout1);


specify
if (B==1'b0 && CI0==1'b1 && CI1==1'b0 && CS==1'b0)
(A => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b0 && CS==1'b1)
(A => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b0)
(A => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b1)
(A => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b0)
(A => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b1)
(A => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b1 && CS==1'b0)
(A => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b1 && CS==1'b1)
(A => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b0 && CS==1'b0)
(B => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b0 && CS==1'b1)
(B => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b0)
(B => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b1)
(B => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b0)
(B => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b1)
(B => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b1 && CS==1'b0)
(B => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b1 && CS==1'b1)
(B => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1==1'b0 && CS==1'b0)
(CI0 => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1==1'b0 && CS==1'b1)
(CI0 => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1==1'b1 && CS==1'b0)
(CI0 => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1==1'b1 && CS==1'b1)
(CI0 => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1==1'b0 && CS==1'b0)
(CI0 => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1==1'b0 && CS==1'b1)
(CI0 => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1==1'b1 && CS==1'b0)
(CI0 => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1==1'b1 && CS==1'b1)
(CI0 => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b0 && CI1==1'b1 && CS==1'b0)
(A => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b0 && CI1==1'b1 && CS==1'b1)
(A => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b0)
(A => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b1)
(A => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b0)
(A => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b1)
(A => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b1 && CI1==1'b0 && CS==1'b0)
(A => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b1 && CI1==1'b0 && CS==1'b1)
(A => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b0 && CI1==1'b1 && CS==1'b0)
(B => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b0 && CI1==1'b1 && CS==1'b1)
(B => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b0)
(B => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b1)
(B => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b0)
(B => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b1)
(B => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b1 && CI1==1'b0 && CS==1'b0)
(B => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b1 && CI1==1'b0 && CS==1'b1)
(B => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0==1'b0 && CS==1'b0)
(CI1 => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0==1'b0 && CS==1'b1)
(CI1 => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0==1'b1 && CS==1'b0)
(CI1 => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0==1'b1 && CS==1'b1)
(CI1 => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0==1'b0 && CS==1'b0)
(CI1 => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0==1'b0 && CS==1'b1)
(CI1 => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0==1'b1 && CS==1'b0)
(CI1 => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0==1'b1 && CS==1'b1)
(CI1 => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b0 && CI1==1'b1 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b0 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b1 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b1 && CI1==1'b0 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b0 && CI1==1'b0 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b0 && CI1==1'b0 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b0 && CI1==1'b1 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b0 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b1 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b1 && CI1==1'b0 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b1 && CI1==1'b1 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b1 && CI1==1'b1 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b0 && CI1==1'b1 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b0 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b1 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b1 && CI1==1'b0 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b0 && CI1==1'b0 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b0 && CI1==1'b0 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b0 && CI1==1'b1 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b0 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b1 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b1 && CI1==1'b0 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b1 && CI1==1'b1 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b1 && CI1==1'b1 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1==1'b0)
(CI0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1==1'b1)
(CI0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1==1'b0)
(CI0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1==1'b1)
(CI0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI1==1'b0)
(CI0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI1==1'b1)
(CI0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI1==1'b0)
(CI0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI1==1'b1)
(CI0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0==1'b0)
(CI1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0==1'b1)
(CI1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0==1'b0)
(CI1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0==1'b1)
(CI1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI0==1'b0)
(CI1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI0==1'b1)
(CI1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI0==1'b0)
(CI1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI0==1'b1)
(CI1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI0==1'b1 && CI1==1'b0)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0==1'b0 && CI1==1'b1)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0==1'b0 && CI1==1'b1)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI0==1'b1 && CI1==1'b0)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI0==1'b0 && CI1==1'b1)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0==1'b1 && CI1==1'b0)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0==1'b1 && CI1==1'b0)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI0==1'b0 && CI1==1'b1)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AFCSHCONX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AFCSHCONX4 (CO0N, CO1N, S, A, B, CI0, CI1, CS);
output S, CO0N, CO1N;
input A, B, CI0, CI1, CS;
  xor I2 (s1, A, B, CI1);
  xor I3 (s2, A, B, CI0);
  and I4 (s3, CS, s1);
  not I5 (csn, CS);
  and I6 (s4, csn, s2);
  or I7 (S, s3, s4);
  and I8 (a_and_b, A, B);
  and I9 (a_and_ci0, A, CI0);
  and I10 (b_and_ci0, B, CI0);
  or I11 (cout0, a_and_b, a_and_ci0, b_and_ci0);
  and I12 (a_and_ci1, A, CI1);
  and I13 (b_and_ci1, B, CI1);
  or I14 (cout1, a_and_b, a_and_ci1, b_and_ci1);
  not I15 (CO0N, cout0);
  not I16 (CO1N, cout1);


specify
if (B==1'b0 && CI0==1'b1 && CI1==1'b0 && CS==1'b0)
(A => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b0 && CS==1'b1)
(A => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b0)
(A => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b1)
(A => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b0)
(A => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b1)
(A => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b1 && CS==1'b0)
(A => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b1 && CS==1'b1)
(A => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b0 && CS==1'b0)
(B => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b0 && CS==1'b1)
(B => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b0)
(B => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b1)
(B => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b0)
(B => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b1)
(B => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b1 && CS==1'b0)
(B => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b1 && CS==1'b1)
(B => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1==1'b0 && CS==1'b0)
(CI0 => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1==1'b0 && CS==1'b1)
(CI0 => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1==1'b1 && CS==1'b0)
(CI0 => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1==1'b1 && CS==1'b1)
(CI0 => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1==1'b0 && CS==1'b0)
(CI0 => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1==1'b0 && CS==1'b1)
(CI0 => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1==1'b1 && CS==1'b0)
(CI0 => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1==1'b1 && CS==1'b1)
(CI0 => CO0N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b0 && CI1==1'b1 && CS==1'b0)
(A => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b0 && CI1==1'b1 && CS==1'b1)
(A => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b0)
(A => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b1)
(A => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b0)
(A => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b1)
(A => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b1 && CI1==1'b0 && CS==1'b0)
(A => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b1 && CI1==1'b0 && CS==1'b1)
(A => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b0 && CI1==1'b1 && CS==1'b0)
(B => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b0 && CI1==1'b1 && CS==1'b1)
(B => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b0)
(B => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b1)
(B => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b0)
(B => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b1)
(B => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b1 && CI1==1'b0 && CS==1'b0)
(B => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b1 && CI1==1'b0 && CS==1'b1)
(B => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0==1'b0 && CS==1'b0)
(CI1 => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0==1'b0 && CS==1'b1)
(CI1 => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0==1'b1 && CS==1'b0)
(CI1 => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0==1'b1 && CS==1'b1)
(CI1 => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0==1'b0 && CS==1'b0)
(CI1 => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0==1'b0 && CS==1'b1)
(CI1 => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0==1'b1 && CS==1'b0)
(CI1 => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0==1'b1 && CS==1'b1)
(CI1 => CO1N) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b0 && CI1==1'b1 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b0 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b1 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b1 && CI1==1'b0 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b0 && CI1==1'b0 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b0 && CI1==1'b0 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b0 && CI1==1'b1 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI0==1'b1 && CI1==1'b0 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b0 && CI1==1'b1 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b1 && CI1==1'b0 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b1 && CI1==1'b1 && CS==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI0==1'b1 && CI1==1'b1 && CS==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b0 && CI1==1'b1 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b0 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b1 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b0 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b1 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b1 && CI1==1'b0 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b0 && CI1==1'b0 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b0 && CI1==1'b0 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b0 && CI1==1'b1 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI0==1'b1 && CI1==1'b0 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b0 && CI1==1'b1 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b1 && CI1==1'b0 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b1 && CI1==1'b1 && CS==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI0==1'b1 && CI1==1'b1 && CS==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1==1'b0)
(CI0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI1==1'b1)
(CI0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1==1'b0)
(CI0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI1==1'b1)
(CI0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI1==1'b0)
(CI0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI1==1'b1)
(CI0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI1==1'b0)
(CI0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI1==1'b1)
(CI0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0==1'b0)
(CI1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0==1'b1)
(CI1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0==1'b0)
(CI1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0==1'b1)
(CI1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI0==1'b0)
(CI1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI0==1'b1)
(CI1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI0==1'b0)
(CI1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI0==1'b1)
(CI1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI0==1'b1 && CI1==1'b0)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0==1'b0 && CI1==1'b1)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0==1'b0 && CI1==1'b1)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI0==1'b1 && CI1==1'b0)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && CI0==1'b0 && CI1==1'b1)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && CI0==1'b1 && CI1==1'b0)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && CI0==1'b1 && CI1==1'b0)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && CI0==1'b0 && CI1==1'b1)
(CS => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AFCSHCONX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AFHCINX2 (CO, S, A, B, CIN);
output S, CO;
input A, B, CIN;
  not I0 (ci, CIN);
  xor I1 (S, A, B, ci);
  and I2 (a_and_b, A, B);
  and I3 (a_and_ci, A, ci);
  and I4 (b_and_ci, B, ci);
  or I5 (CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CIN==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CIN==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CIN==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CIN => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CIN => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CIN => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CIN => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AFHCINX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AFHCINX4 (CO, S, A, B, CIN);
output S, CO;
input A, B, CIN;
  not I0 (ci, CIN);
  xor I1 (S, A, B, ci);
  and I2 (a_and_b, A, B);
  and I3 (a_and_ci, A, ci);
  and I4 (b_and_ci, B, ci);
  or I5 (CO, a_and_b, a_and_ci, b_and_ci);


specify
if (B==1'b0 && CIN==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CIN==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CIN==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CIN==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CIN==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CIN==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CIN => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CIN => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CIN => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CIN => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AFHCINX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AFHCONX2 (CON, S, A, B, CI);
output S, CON;
input A, B, CI;
  xor I0 (S, A, B, CI);
  and I1 (a_and_b, A, B);
  and I2 (a_and_ci, A, CI);
  and I3 (b_and_ci, B, CI);
  or I4 (cout, a_and_b, a_and_ci, b_and_ci);
  not I5 (CON, cout);


specify
if (B==1'b0 && CI==1'b1)
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AFHCONX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AFHCONX4 (CON, S, A, B, CI);
output S, CON;
input A, B, CI;
  xor I0 (S, A, B, CI);
  and I1 (a_and_b, A, B);
  and I2 (a_and_ci, A, CI);
  and I3 (b_and_ci, B, CI);
  or I4 (cout, a_and_b, a_and_ci, b_and_ci);
  not I5 (CON, cout);


specify
if (B==1'b0 && CI==1'b1)
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && CI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && CI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && CI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && CI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(CI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AFHCONX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AHHCINX2 (CO, S, A, CIN);
output S, CO;
input A, CIN;
  not I0 (ci, CIN);
  xor I1 (S, A, ci);
  and I2 (CO, A, ci);


specify
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CIN => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge CIN => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AHHCINX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AHHCINX4 (CO, S, A, CIN);
output S, CO;
input A, CIN;
  not I0 (ci, CIN);
  xor I1 (S, A, ci);
  and I2 (CO, A, ci);


specify
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(CIN => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CIN => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge CIN => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AHHCINX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AHHCONX2 (CON, S, A, CI);
output S, CON;
input A, CI;
  xor I0 (S, A, CI);
  and  I1 (cout, A, CI);
  not I2 (CON, cout);


specify
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CI => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge CI => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AHHCONX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AHHCONX4 (CON, S, A, CI);
output S, CON;
input A, CI;
  xor I0 (S, A, CI);
  and  I1 (cout, A, CI);
  not I2 (CON, cout);


specify
(A => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(CI => CON) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CI => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge CI => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AHHCONX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2X1 (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2X2 (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2X4 (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND2XL (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND2XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3X1 (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3X2 (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3X4 (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND3XL (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND3XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4X1 (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4X2 (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4X4 (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AND4XL (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AND4XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module ANTENNA (A);
input A;

specify

endspecify
endmodule // ANTENNA
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211X1 (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI211X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211X2 (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI211X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211X4 (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI211X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI211XL (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI211XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21X1 (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21X2 (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21X4 (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI21XL (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI21XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221X1 (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, C0, outB, outA);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI221X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221X2 (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, C0, outB, outA);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI221X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221X4 (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, C0, outB, outA);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI221X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI221XL (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, C0, outB, outA);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI221XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222X1 (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(Y, outA, outB, outC);


specify
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI222X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222X2 (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(Y, outA, outB, outC);


specify
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI222X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222X4 (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(Y, outA, outB, outC);


specify
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI222X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI222XL (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(Y, outA, outB, outC);


specify
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI222XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22X1 (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22X2 (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22X4 (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI22XL (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI22XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB1X1 (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;



  nor I0 (outA, A0N, A1N);
  nor I1 (Y, B0, outA);


specify
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB1X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB1X2 (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;



  nor I0 (outA, A0N, A1N);
  nor I1 (Y, B0, outA);


specify
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB1X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB1X4 (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;



  nor I0 (outA, A0N, A1N);
  nor I1 (Y, B0, outA);


specify
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB1X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB1XL (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;



  nor I0 (outA, A0N, A1N);
  nor I1 (Y, B0, outA);


specify
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB1XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB2X1 (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;



  nor I0 (outA, A0N, A1N);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB2X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB2X2 (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;



  nor I0 (outA, A0N, A1N);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB2X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB2X4 (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;



  nor I0 (outA, A0N, A1N);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB2X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI2BB2XL (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;



  nor I0 (outA, A0N, A1N);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI2BB2XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31X1 (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI31X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31X2 (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI31X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31X4 (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI31X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI31XL (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  and I0(outA, A0, A1, A2);
  nor I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI31XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32X1 (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI32X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32X2 (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI32X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32X4 (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI32X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI32XL (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI32XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI33X1 (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1, B2);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI33X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI33X2 (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1, B2);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI33X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI33X4 (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1, B2);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI33X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module AOI33XL (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;



  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1, B2);
  nor I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // AOI33XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BENCX1 (A, S, X2, M0, M1, M2);
output S, A, X2;
input M2, M1, M0;

  not I0 (m1n, M1);
  not I1 (m0n, M0);
  or  I3 (m1n_or_m0n, m1n, m0n);
  nand I4 (S, M2, m1n_or_m0n);
  or  I5 (m1_or_m0, M1, M0);
  nand I6 (A, m2n, m1_or_m0);
  xor I7 (x2n, M1, M0);
  not I8 (X2, x2n);
  not I9 (m2n, M2);



specify
(M0 => A) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => A) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => A) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => A) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b1)
(M2 => A) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b0)
(M2 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BENCX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BENCX2 (A, S, X2, M0, M1, M2);
output S, A, X2;
input M2, M1, M0;

  not I0 (m1n, M1);
  not I1 (m0n, M0);
  or  I3 (m1n_or_m0n, m1n, m0n);
  nand I4 (S, M2, m1n_or_m0n);
  or  I5 (m1_or_m0, M1, M0);
  nand I6 (A, m2n, m1_or_m0);
  xor I7 (x2n, M1, M0);
  not I8 (X2, x2n);
  not I9 (m2n, M2);



specify
(M0 => A) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => A) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => A) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => A) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b1)
(M2 => A) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b0)
(M2 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BENCX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BENCX4 (A, S, X2, M0, M1, M2);
output S, A, X2;
input M2, M1, M0;

  not I0 (m1n, M1);
  not I1 (m0n, M0);
  or  I3 (m1n_or_m0n, m1n, m0n);
  nand I4 (S, M2, m1n_or_m0n);
  or  I5 (m1_or_m0, M1, M0);
  nand I6 (A, m2n, m1_or_m0);
  xor I7 (x2n, M1, M0);
  not I8 (X2, x2n);
  not I9 (m2n, M2);



specify
(M0 => A) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => A) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => A) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => A) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b1)
(M2 => A) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M0 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(M1 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b0)
(M2 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1)
(M2 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0)
(M2 => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M0 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b0)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(posedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M2==1'b1)
(negedge M1 => (X2:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BENCX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BMXX1 (PP, A, M0, M1, S, X2);
output PP;
input X2, A, S, M1, M0;

  udp_bmx I0 (PP, X2, A, S, M1, M0);



specify
if (M0==1'b0 && M1==1'b1 && S==1'b0 && X2==1'b0)
(A => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0 && M1==1'b1 && S==1'b1 && X2==1'b0)
(A => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0 && S==1'b0 && X2==1'b1)
(A => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b0 && S==1'b1 && X2==1'b1)
(A => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b1 && S==1'b0 && X2==1'b0)
(A => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b1 && S==1'b0 && X2==1'b1)
(A => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b1 && S==1'b1 && X2==1'b0)
(A => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1 && M1==1'b1 && S==1'b1 && X2==1'b1)
(A => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M1==1'b0)
(posedge M0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M1==1'b0)
(negedge M0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M1==1'b1)
(posedge M0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M1==1'b1)
(negedge M0 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0)
(posedge M1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b0)
(negedge M1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1)
(posedge M1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (M0==1'b1)
(negedge M1 => (PP:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && M0==1'b0 && M1==1'b0 && X2==1'b0)
(S => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && M0==1'b0 && M1==1'b0 && X2==1'b1)
(S => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && M0==1'b0 && M1==1'b1 && X2==1'b1)
(S => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && M0==1'b1 && M1==1'b0 && X2==1'b0)
(S => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && M0==1'b0 && M1==1'b0 && X2==1'b0)
(S => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && M0==1'b0 && M1==1'b0 && X2==1'b1)
(S => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && M0==1'b0 && M1==1'b1 && X2==1'b1)
(S => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && M0==1'b1 && M1==1'b0 && X2==1'b0)
(S => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && M0==1'b0 && M1==1'b1 && S==1'b1)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && M0==1'b1 && M1==1'b0 && S==1'b0)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && M0==1'b1 && M1==1'b0 && S==1'b1)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && M0==1'b0 && M1==1'b1 && S==1'b0)
(X2 => PP) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BMXX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFX1 (Y, A);
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFX12 (Y, A);
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFX12
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFX16 (Y, A);
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFX16
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFX2 (Y, A);
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFX20 (Y, A);
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFX20
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFX3 (Y, A);
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFX3
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFX4 (Y, A);
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFX8 (Y, A);
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFX8
`endcelldefine
`timescale 1ns/1ps
`celldefine
module BUFXL (Y, A);
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // BUFXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUFX1 (Y, A);
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUFX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUFX12 (Y, A);
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUFX12
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUFX16 (Y, A);
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUFX16
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUFX2 (Y, A);
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUFX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUFX20 (Y, A);
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUFX20
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUFX3 (Y, A);
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUFX3
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUFX4 (Y, A);
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUFX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUFX8 (Y, A);
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUFX8
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKBUFXL (Y, A);
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKBUFXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINVX1 (Y, A);
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINVX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINVX12 (Y, A);
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINVX12
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINVX16 (Y, A);
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINVX16
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINVX2 (Y, A);
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINVX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINVX20 (Y, A);
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINVX20
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINVX3 (Y, A);
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINVX3
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINVX4 (Y, A);
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINVX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINVX8 (Y, A);
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINVX8
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CLKINVXL (Y, A);
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CLKINVXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CMPR22X1 (CO, S, A, B);
output S, CO;
input A, B;
  xor I0(S, A, B);
  and I1(CO, A, B);


specify
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (S:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CMPR22X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CMPR32X1 (CO, S, A, B, C);
output S, CO;
input A, B, C;

  xor I0 (t1, A, B);
  xor I1 (S, t1, C);
  and I2 (t2, A, B);
  and I3 (t3, t1, C);
  or  I4 (CO, t2, t3);



specify
if (B==1'b0 && C==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CMPR32X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CMPR42X1 (CO, ICO, S, A, B, C, D, ICI);
output S, CO, ICO;
input A, B, C, D, ICI;

  xor I0 (t1, A, B);
  xor I1 (IS, t1, C);
  and I2 (t2, A, B);
  and I3 (t3, A, C);
  and I4 (t4, B, C);
  or   I5 (ICO, t2, t3, t4);
  xor I6 (ss, IS, D);
  xor  I7 (S, ss, ICI);
  and I8 (t5, IS, D);
  and I9 (t6, IS, ICI);
  and I10 (t7, D, ICI);
  or   I11 (CO, t5, t6, t7);



specify
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0 && ICI==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1 && ICI==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0 && ICI==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1 && ICI==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && ICI==1'b1)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && ICI==1'b0)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && ICI==1'b0)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && ICI==1'b1)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && ICI==1'b0)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && ICI==1'b1)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && ICI==1'b1)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && ICI==1'b0)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && ICI==1'b0)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && ICI==1'b1)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && ICI==1'b1)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && ICI==1'b0)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && ICI==1'b1)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && ICI==1'b0)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && ICI==1'b0)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && ICI==1'b1)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b0)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b1)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CMPR42X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module CMPR42X2 (CO, ICO, S, A, B, C, D, ICI);
output S, CO, ICO;
input A, B, C, D, ICI;

  xor I0 (t1, A, B);
  xor I1 (IS, t1, C);
  and I2 (t2, A, B);
  and I3 (t3, A, C);
  and I4 (t4, B, C);
  or   I5 (ICO, t2, t3, t4);
  xor I6 (ss, IS, D);
  xor  I7 (S, ss, ICI);
  and I8 (t5, IS, D);
  and I9 (t6, IS, ICI);
  and I10 (t7, D, ICI);
  or   I11 (CO, t5, t6, t7);



specify
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && ICI==1'b1)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && ICI==1'b0)
(D => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0)
(ICI => CO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(A => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(B => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b1)
(C => ICO) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b0)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b1)
(A => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0 && ICI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1 && ICI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0 && ICI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1 && ICI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0 && ICI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1 && ICI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0 && ICI==1'b0)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1 && ICI==1'b1)
(B => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0 && ICI==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1 && ICI==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0 && ICI==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1 && ICI==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0 && ICI==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1 && ICI==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0 && ICI==1'b0)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1 && ICI==1'b1)
(C => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && ICI==1'b1)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && ICI==1'b0)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && ICI==1'b0)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && ICI==1'b1)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && ICI==1'b0)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && ICI==1'b1)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && ICI==1'b1)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && ICI==1'b0)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && ICI==1'b0)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && ICI==1'b1)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && ICI==1'b1)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && ICI==1'b0)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && ICI==1'b1)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && ICI==1'b0)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && ICI==1'b0)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && ICI==1'b1)
(D => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b0)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b1)
(ICI => S) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // CMPR42X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DFFHQX1 (Q, CK, D);
output Q;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);


specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFHQX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFHQX2 (Q, CK, D);
output Q;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);


specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFHQX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFHQX4 (Q, CK, D);
output Q;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);


specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFHQX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFHQXL (Q, CK, D);
output Q;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);


specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFHQXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNRX1 (Q, QN, CKN, D, RN);
output Q, QN;
input  D, CKN, RN;
reg NOTIFIER;
supply1 xSN;

  buf   XX0 (xRN, RN);
  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_D ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, negedge CKN &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // DFFNRX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNRX2 (Q, QN, CKN, D, RN);
output Q, QN;
input  D, CKN, RN;
reg NOTIFIER;
supply1 xSN;

  buf   XX0 (xRN, RN);
  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_D ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, negedge CKN &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // DFFNRX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNRX4 (Q, QN, CKN, D, RN);
output Q, QN;
input  D, CKN, RN;
reg NOTIFIER;
supply1 xSN;

  buf   XX0 (xRN, RN);
  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_D ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, negedge CKN &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // DFFNRX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNRXL (Q, QN, CKN, D, RN);
output Q, QN;
input  D, CKN, RN;
reg NOTIFIER;
supply1 xSN;

  buf   XX0 (xRN, RN);
  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_D ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, negedge CKN &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // DFFNRXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSRX1 (Q, QN, CKN, D, RN, SN);
output Q, QN;
input  D, CKN, SN, RN;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  not      IC (clk, CKN);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, negedge CKN &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFNSRX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSRX2 (Q, QN, CKN, D, RN, SN);
output Q, QN;
input  D, CKN, SN, RN;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  not      IC (clk, CKN);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, negedge CKN &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFNSRX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSRX4 (Q, QN, CKN, D, RN, SN);
output Q, QN;
input  D, CKN, SN, RN;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  not      IC (clk, CKN);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, negedge CKN &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFNSRX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSRXL (Q, QN, CKN, D, RN, SN);
output Q, QN;
input  D, CKN, SN, RN;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  not      IC (clk, CKN);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, negedge CKN &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFNSRXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSX1 (Q, QN, CKN, D, SN);
output Q, QN;
input  D, CKN, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFNSX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSX2 (Q, QN, CKN, D, SN);
output Q, QN;
input  D, CKN, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFNSX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSX4 (Q, QN, CKN, D, SN);
output Q, QN;
input  D, CKN, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFNSX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNSXL (Q, QN, CKN, D, SN);
output Q, QN;
input  D, CKN, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFNSXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNX1 (Q, QN, CKN, D);
output Q, QN;
input  D, CKN;
reg NOTIFIER;
supply1 xSN,xRN;
  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);


specify
$width(posedge CKN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFNX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNX2 (Q, QN, CKN, D);
output Q, QN;
input  D, CKN;
reg NOTIFIER;
supply1 xSN,xRN;
  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);


specify
$width(posedge CKN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFNX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNX4 (Q, QN, CKN, D);
output Q, QN;
input  D, CKN;
reg NOTIFIER;
supply1 xSN,xRN;
  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);


specify
$width(posedge CKN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFNX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFNXL (Q, QN, CKN, D);
output Q, QN;
input  D, CKN;
reg NOTIFIER;
supply1 xSN,xRN;
  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);


specify
$width(posedge CKN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(negedge CKN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge CKN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFNXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRHQX1 (Q, CK, D, RN);
output Q;
input  D, CK, RN;
reg NOTIFIER;
supply1 xSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_RN ;
wire ENABLE_D ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFRHQX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRHQX2 (Q, CK, D, RN);
output Q;
input  D, CK, RN;
reg NOTIFIER;
supply1 xSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_RN ;
wire ENABLE_D ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFRHQX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRHQX4 (Q, CK, D, RN);
output Q;
input  D, CK, RN;
reg NOTIFIER;
supply1 xSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_RN ;
wire ENABLE_D ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFRHQX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRHQXL (Q, CK, D, RN);
output Q;
input  D, CK, RN;
reg NOTIFIER;
supply1 xSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_RN ;
wire ENABLE_D ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFRHQXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRX1 (Q, QN, CK, D, RN);
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
supply1 xSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_D ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // DFFRX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRX2 (Q, QN, CK, D, RN);
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
supply1 xSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_D ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // DFFRX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRX4 (Q, QN, CK, D, RN);
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
supply1 xSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_D ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // DFFRX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFRXL (Q, QN, CK, D, RN);
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
supply1 xSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_D ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // DFFRXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSHQX1 (Q, CK, D, SN);
output Q;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // DFFSHQX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSHQX2 (Q, CK, D, SN);
output Q;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // DFFSHQX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSHQX4 (Q, CK, D, SN);
output Q;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // DFFSHQX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSHQXL (Q, CK, D, SN);
output Q;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // DFFSHQXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRHQX1 (Q, CK, D, RN, SN);
output Q;
input  D, CK, SN, RN;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // DFFSRHQX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRHQX2 (Q, CK, D, RN, SN);
output Q;
input  D, CK, SN, RN;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // DFFSRHQX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRHQX4 (Q, CK, D, RN, SN);
output Q;
input  D, CK, SN, RN;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // DFFSRHQX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRHQXL (Q, CK, D, RN, SN);
output Q;
input  D, CK, SN, RN;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // DFFSRHQXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRX1 (Q, QN, CK, D, RN, SN);
output Q, QN;
input  D, CK, SN, RN;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSRX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRX2 (Q, QN, CK, D, RN, SN);
output Q, QN;
input  D, CK, SN, RN;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSRX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRX4 (Q, QN, CK, D, RN, SN);
output Q, QN;
input  D, CK, SN, RN;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSRX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSRXL (Q, QN, CK, D, RN, SN);
output Q, QN;
input  D, CK, SN, RN;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  buf   XX1 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSRXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSX1 (Q, QN, CK, D, SN);
output Q, QN;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSX2 (Q, QN, CK, D, SN);
output Q, QN;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSX4 (Q, QN, CK, D, SN);
output Q, QN;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFSXL (Q, QN, CK, D, SN);
output Q, QN;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // DFFSXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFTRX1 (Q, QN, CK, D, RN);
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
supply1 xSN, EN,flag;

  buf   XX0 (xRN, RN);
  and F0 (rn_and_sn, xRN,xSN);
  buf     IC (clk, CK);
  udp_edfft I0 (n0, D, clk, xRN, xSN, EN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_D ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (RN==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (RN==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFTRX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFTRX2 (Q, QN, CK, D, RN);
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
supply1 xSN, EN,flag;

  buf   XX0 (xRN, RN);
  and F0 (rn_and_sn, xRN,xSN);
  buf     IC (clk, CK);
  udp_edfft I0 (n0, D, clk, xRN, xSN, EN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_D ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (RN==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (RN==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFTRX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFTRX4 (Q, QN, CK, D, RN);
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
supply1 xSN, EN,flag;

  buf   XX0 (xRN, RN);
  and F0 (rn_and_sn, xRN,xSN);
  buf     IC (clk, CK);
  udp_edfft I0 (n0, D, clk, xRN, xSN, EN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_D ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (RN==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (RN==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFTRX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFTRXL (Q, QN, CK, D, RN);
output Q, QN;
input  D, CK, RN;
reg NOTIFIER;
supply1 xSN, EN,flag;

  buf   XX0 (xRN, RN);
  and F0 (rn_and_sn, xRN,xSN);
  buf     IC (clk, CK);
  udp_edfft I0 (n0, D, clk, xRN, xSN, EN, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_D ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (RN==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (RN==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFTRXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFX1 (Q, QN, CK, D);
output Q, QN;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);


specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFX1
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFX2 (Q, QN, CK, D);
output Q, QN;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);


specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFX2
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFX4 (Q, QN, CK, D);
output Q, QN;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);


specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFX4
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DFFXL (Q, QN, CK, D);
output Q, QN;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);


specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DFFXL
`endcelldefine

`timescale 1ns/1ps
`celldefine
module DLY1X1 (Y, A);
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLY1X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLY2X1 (Y, A);
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLY2X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLY3X1 (Y, A);
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLY3X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module DLY4X1 (Y, A);
output Y;
input A;

  buf I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // DLY4X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module EDFFTRX1 (Q, QN, CK, D, E, RN);
output Q, QN;
input D, CK, E, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

  udp_edfft I0 (n0, D, CK, xRN, xSN, E, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_E_OR_NOT_RN ;
wire ENABLE_E_AND_RN ;
wire ENABLE_RN ;
wire ENABLE_D_OR_NOT_E ;
assign ENABLE_E_OR_NOT_RN = (E | !RN) ? 1'b1:1'b0;
assign ENABLE_E_AND_RN = (E&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D_OR_NOT_E = (D | !E) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_NOT_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_NOT_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_OR_NOT_E == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_OR_NOT_E == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (E==1'b1 && RN==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFFTRX1
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFFTRX2 (Q, QN, CK, D, E, RN);
output Q, QN;
input D, CK, E, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

  udp_edfft I0 (n0, D, CK, xRN, xSN, E, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_E_OR_NOT_RN ;
wire ENABLE_E_AND_RN ;
wire ENABLE_RN ;
wire ENABLE_D_OR_NOT_E ;
assign ENABLE_E_OR_NOT_RN = (E | !RN) ? 1'b1:1'b0;
assign ENABLE_E_AND_RN = (E&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D_OR_NOT_E = (D | !E) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_NOT_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_NOT_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_OR_NOT_E == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_OR_NOT_E == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (E==1'b1 && RN==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFFTRX2
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFFTRX4 (Q, QN, CK, D, E, RN);
output Q, QN;
input D, CK, E, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

  udp_edfft I0 (n0, D, CK, xRN, xSN, E, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_E_OR_NOT_RN ;
wire ENABLE_E_AND_RN ;
wire ENABLE_RN ;
wire ENABLE_D_OR_NOT_E ;
assign ENABLE_E_OR_NOT_RN = (E | !RN) ? 1'b1:1'b0;
assign ENABLE_E_AND_RN = (E&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D_OR_NOT_E = (D | !E) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_NOT_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_NOT_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_OR_NOT_E == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_OR_NOT_E == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (E==1'b1 && RN==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFFTRX4
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFFTRXL (Q, QN, CK, D, E, RN);
output Q, QN;
input D, CK, E, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

  udp_edfft I0 (n0, D, CK, xRN, xSN, E, NOTIFIER);
  buf     I1 (Q, n0);
  not     I2 (QN, n0);

wire ENABLE_E_OR_NOT_RN ;
wire ENABLE_E_AND_RN ;
wire ENABLE_RN ;
wire ENABLE_D_OR_NOT_E ;
assign ENABLE_E_OR_NOT_RN = (E | !RN) ? 1'b1:1'b0;
assign ENABLE_E_AND_RN = (E&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D_OR_NOT_E = (D | !E) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_NOT_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_NOT_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_OR_NOT_E == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_OR_NOT_E == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (E==1'b1 && RN==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFFTRXL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFFX1 (Q, QN, CK, D, E);
output Q, QN;
input D, CK, E;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff_PWR I0 (n0, D, CK, xRN, xSN, E, 1'b1, 1'b0, NOTIFIER);
  buf     B1 (Q, n0);
  not      I1 (QN, n0);

wire ENABLE_E ;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFFX1
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFFX2 (Q, QN, CK, D, E);
output Q, QN;
input D, CK, E;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff_PWR I0 (n0, D, CK, xRN, xSN, E, 1'b1, 1'b0, NOTIFIER);
  buf     B1 (Q, n0);
  not      I1 (QN, n0);

wire ENABLE_E ;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFFX2
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFFX4 (Q, QN, CK, D, E);
output Q, QN;
input D, CK, E;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff_PWR I0 (n0, D, CK, xRN, xSN, E, 1'b1, 1'b0, NOTIFIER);
  buf     B1 (Q, n0);
  not      I1 (QN, n0);

wire ENABLE_E ;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFFX4
`endcelldefine


`timescale 1ns/1ps
`celldefine
module EDFFXL (Q, QN, CK, D, E);
output Q, QN;
input D, CK, E;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff_PWR I0 (n0, D, CK, xRN, xSN, E, 1'b1, 1'b0, NOTIFIER);
  buf     B1 (Q, n0);
  not      I1 (QN, n0);

wire ENABLE_E ;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // EDFFXL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module FILL1;
endmodule //FILL1

`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILL16;
endmodule //FILL16

`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILL2;
endmodule //FILL2

`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILL32;
endmodule //FILL32

`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILL4;
endmodule //FILL4

`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILL64;
endmodule //FILL64

`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILL8;
endmodule //FILL8

`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILLCAP16;

specify

endspecify
endmodule // FILLCAP16
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILLCAP3;

specify

endspecify
endmodule // FILLCAP3
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILLCAP32;

specify

endspecify
endmodule // FILLCAP32
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILLCAP4;

specify

endspecify
endmodule // FILLCAP4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILLCAP5;

specify

endspecify
endmodule // FILLCAP5
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILLCAP64;

specify

endspecify
endmodule // FILLCAP64
`endcelldefine
`timescale 1ns/1ps
`celldefine
module FILLCAP8;

specify

endspecify
endmodule // FILLCAP8
`endcelldefine
`timescale 1ns/1ps
`celldefine
module HOLDX1 (Y);
inout Y;

wire io_wire;

  buf(weak0,weak1) I0(Y, io_wire);
  buf I1(io_wire, Y);



specify

endspecify
endmodule // HOLDX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INVX1 (Y, A);
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INVX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INVX12 (Y, A);
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INVX12
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INVX16 (Y, A);
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INVX16
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INVX2 (Y, A);
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INVX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INVX20 (Y, A);
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INVX20
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INVX3 (Y, A);
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INVX3
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INVX4 (Y, A);
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INVX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INVX8 (Y, A);
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INVX8
`endcelldefine
`timescale 1ns/1ps
`celldefine
module INVXL (Y, A);
output Y;
input A;

  not I0(Y, A);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // INVXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module JKFFRX1 (Q, QN, CK, J, K, RN);
output Q, QN;
input  J, K, CK, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);

udp_jkff_PWR I0 (n0,J, K,CK, xRN, xSN, 1'b1, 1'b0, NOTIFIER); 
buf I1 (Q,n0);
not I2 (QN,n0);

wire ENABLE_J_AND_RN_OR_K_AND_RN ;
wire ENABLE_RN ;
wire ENABLE_J ;
assign ENABLE_J_AND_RN_OR_K_AND_RN = (J&RN | K&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_J = (J) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_J_AND_RN_OR_K_AND_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_J_AND_RN_OR_K_AND_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_J == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // JKFFRX1
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFRX2 (Q, QN, CK, J, K, RN);
output Q, QN;
input  J, K, CK, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);

udp_jkff_PWR I0 (n0,J, K,CK, xRN, xSN, 1'b1, 1'b0, NOTIFIER); 
buf I1 (Q,n0);
not I2 (QN,n0);

wire ENABLE_J_AND_RN_OR_K_AND_RN ;
wire ENABLE_RN ;
wire ENABLE_J ;
assign ENABLE_J_AND_RN_OR_K_AND_RN = (J&RN | K&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_J = (J) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_J_AND_RN_OR_K_AND_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_J_AND_RN_OR_K_AND_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_J == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // JKFFRX2
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFRX4 (Q, QN, CK, J, K, RN);
output Q, QN;
input  J, K, CK, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);

udp_jkff_PWR I0 (n0,J, K,CK, xRN, xSN, 1'b1, 1'b0, NOTIFIER); 
buf I1 (Q,n0);
not I2 (QN,n0);

wire ENABLE_J_AND_RN_OR_K_AND_RN ;
wire ENABLE_RN ;
wire ENABLE_J ;
assign ENABLE_J_AND_RN_OR_K_AND_RN = (J&RN | K&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_J = (J) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_J_AND_RN_OR_K_AND_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_J_AND_RN_OR_K_AND_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_J == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // JKFFRX4
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFRXL (Q, QN, CK, J, K, RN);
output Q, QN;
input  J, K, CK, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);

udp_jkff_PWR I0 (n0,J, K,CK, xRN, xSN, 1'b1, 1'b0, NOTIFIER); 
buf I1 (Q,n0);
not I2 (QN,n0);

wire ENABLE_J_AND_RN_OR_K_AND_RN ;
wire ENABLE_RN ;
wire ENABLE_J ;
assign ENABLE_J_AND_RN_OR_K_AND_RN = (J&RN | K&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_J = (J) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_J_AND_RN_OR_K_AND_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_J_AND_RN_OR_K_AND_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), posedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN == 1'b1), negedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_J == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // JKFFRXL
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFSRX1 (Q, QN, CK, J, K, RN, SN);
output Q, QN;
input  J, K, CK, SN, RN;
reg NOTIFIER;

  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);

udp_jkff I0 (n0,J, K,CK, xRN, xSN, NOTIFIER); 
buf I1 (Q,n0);
not I2 (QN,n0);

wire ENABLE_J_AND_RN_AND_SN_OR_K_AND_RN_AND_SN ;
wire ENABLE_RN_AND_SN ;
wire ENABLE_J_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_K_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_J_AND_RN_AND_SN_OR_K_AND_RN_AND_SN = (J&RN&SN | K&RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_J_AND_SN = (J&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_K_AND_RN = (K&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_J_AND_RN_AND_SN_OR_K_AND_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_J_AND_RN_AND_SN_OR_K_AND_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_J_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_K_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // JKFFSRX1
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFSRX2 (Q, QN, CK, J, K, RN, SN);
output Q, QN;
input  J, K, CK, SN, RN;
reg NOTIFIER;

  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);

udp_jkff I0 (n0,J, K,CK, xRN, xSN, NOTIFIER); 
buf I1 (Q,n0);
not I2 (QN,n0);

wire ENABLE_J_AND_RN_AND_SN_OR_K_AND_RN_AND_SN ;
wire ENABLE_RN_AND_SN ;
wire ENABLE_J_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_K_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_J_AND_RN_AND_SN_OR_K_AND_RN_AND_SN = (J&RN&SN | K&RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_J_AND_SN = (J&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_K_AND_RN = (K&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_J_AND_RN_AND_SN_OR_K_AND_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_J_AND_RN_AND_SN_OR_K_AND_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_J_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_K_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // JKFFSRX2
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFSRX4 (Q, QN, CK, J, K, RN, SN);
output Q, QN;
input  J, K, CK, SN, RN;
reg NOTIFIER;

  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);

udp_jkff I0 (n0,J, K,CK, xRN, xSN, NOTIFIER); 
buf I1 (Q,n0);
not I2 (QN,n0);

wire ENABLE_J_AND_RN_AND_SN_OR_K_AND_RN_AND_SN ;
wire ENABLE_RN_AND_SN ;
wire ENABLE_J_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_K_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_J_AND_RN_AND_SN_OR_K_AND_RN_AND_SN = (J&RN&SN | K&RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_J_AND_SN = (J&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_K_AND_RN = (K&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_J_AND_RN_AND_SN_OR_K_AND_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_J_AND_RN_AND_SN_OR_K_AND_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_J_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_K_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // JKFFSRX4
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFSRXL (Q, QN, CK, J, K, RN, SN);
output Q, QN;
input  J, K, CK, SN, RN;
reg NOTIFIER;

  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);

udp_jkff I0 (n0,J, K,CK, xRN, xSN, NOTIFIER); 
buf I1 (Q,n0);
not I2 (QN,n0);

wire ENABLE_J_AND_RN_AND_SN_OR_K_AND_RN_AND_SN ;
wire ENABLE_RN_AND_SN ;
wire ENABLE_J_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_K_AND_RN ;
wire ENABLE_RN ;
assign ENABLE_J_AND_RN_AND_SN_OR_K_AND_RN_AND_SN = (J&RN&SN | K&RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_J_AND_SN = (J&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_K_AND_RN = (K&RN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_J_AND_RN_AND_SN_OR_K_AND_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_J_AND_RN_AND_SN_OR_K_AND_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), posedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), negedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_J_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_K_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // JKFFSRXL
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFSX1 (Q, QN, CK, J, K, SN);
output Q, QN;
input  J, K, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;
  buf   XX0 (xSN, SN);

udp_jkff_PWR I0 (n0,J, K,CK, xRN, xSN, 1'b1, 1'b0, NOTIFIER); 
buf I1 (Q,n0);
not I2 (QN,n0);

wire ENABLE_J_AND_SN_OR_K_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_K ;
assign ENABLE_J_AND_SN_OR_K_AND_SN = (J&SN | K&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_K = (K) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_J_AND_SN_OR_K_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_J_AND_SN_OR_K_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_K == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // JKFFSX1
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFSX2 (Q, QN, CK, J, K, SN);
output Q, QN;
input  J, K, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;
  buf   XX0 (xSN, SN);

udp_jkff_PWR I0 (n0,J, K,CK, xRN, xSN, 1'b1, 1'b0, NOTIFIER); 
buf I1 (Q,n0);
not I2 (QN,n0);

wire ENABLE_J_AND_SN_OR_K_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_K ;
assign ENABLE_J_AND_SN_OR_K_AND_SN = (J&SN | K&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_K = (K) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_J_AND_SN_OR_K_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_J_AND_SN_OR_K_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_K == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // JKFFSX2
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFSX4 (Q, QN, CK, J, K, SN);
output Q, QN;
input  J, K, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;
  buf   XX0 (xSN, SN);

udp_jkff_PWR I0 (n0,J, K,CK, xRN, xSN, 1'b1, 1'b0, NOTIFIER); 
buf I1 (Q,n0);
not I2 (QN,n0);

wire ENABLE_J_AND_SN_OR_K_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_K ;
assign ENABLE_J_AND_SN_OR_K_AND_SN = (J&SN | K&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_K = (K) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_J_AND_SN_OR_K_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_J_AND_SN_OR_K_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_K == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // JKFFSX4
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFSXL (Q, QN, CK, J, K, SN);
output Q, QN;
input  J, K, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;
  buf   XX0 (xSN, SN);

udp_jkff_PWR I0 (n0,J, K,CK, xRN, xSN, 1'b1, 1'b0, NOTIFIER); 
buf I1 (Q,n0);
not I2 (QN,n0);

wire ENABLE_J_AND_SN_OR_K_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_K ;
assign ENABLE_J_AND_SN_OR_K_AND_SN = (J&SN | K&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_K = (K) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_J_AND_SN_OR_K_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_J_AND_SN_OR_K_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), posedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SN == 1'b1), negedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_K == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b0 && K==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && J==1'b1 && K==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b0 && K==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && J==1'b1 && K==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // JKFFSXL
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFX1 (Q, QN, CK, J, K);
output Q, QN;
input  J, K, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

udp_jkff_PWR I0 (n0,J, K,CK, xRN, xSN, 1'b1, 1'b0, NOTIFIER); 
buf I1 (Q,n0);
not I2 (QN,n0);

wire ENABLE_J_OR_K ;
assign ENABLE_J_OR_K = (J | K) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_J_OR_K == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_J_OR_K == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, posedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // JKFFX1
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFX2 (Q, QN, CK, J, K);
output Q, QN;
input  J, K, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

udp_jkff_PWR I0 (n0,J, K,CK, xRN, xSN, 1'b1, 1'b0, NOTIFIER); 
buf I1 (Q,n0);
not I2 (QN,n0);

wire ENABLE_J_OR_K ;
assign ENABLE_J_OR_K = (J | K) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_J_OR_K == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_J_OR_K == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, posedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // JKFFX2
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFX4 (Q, QN, CK, J, K);
output Q, QN;
input  J, K, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

udp_jkff_PWR I0 (n0,J, K,CK, xRN, xSN, 1'b1, 1'b0, NOTIFIER); 
buf I1 (Q,n0);
not I2 (QN,n0);

wire ENABLE_J_OR_K ;
assign ENABLE_J_OR_K = (J | K) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_J_OR_K == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_J_OR_K == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, posedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // JKFFX4
`endcelldefine





`timescale 1ns/1ps
`celldefine
module JKFFXL (Q, QN, CK, J, K);
output Q, QN;
input  J, K, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

udp_jkff_PWR I0 (n0,J, K,CK, xRN, xSN, 1'b1, 1'b0, NOTIFIER); 
buf I1 (Q,n0);
not I2 (QN,n0);

wire ENABLE_J_OR_K ;
assign ENABLE_J_OR_K = (J | K) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_J_OR_K == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_J_OR_K == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge J, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, posedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge K, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b0 || J==1'b0 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (J==1'b1 && K==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // JKFFXL
`endcelldefine





`timescale 1ns/1ps
`celldefine
module MX2X1 (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2X2 (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2X4 (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX2XL (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX2XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX4X1 (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(Y, A, B, C, D, S0, S1);



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX4X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX4X2 (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(Y, A, B, C, D, S0, S1);



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX4X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX4X4 (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(Y, A, B, C, D, S0, S1);



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX4X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MX4XL (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(Y, A, B, C, D, S0, S1);



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MX4XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2X1 (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI2X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2X2 (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI2X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2X4 (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI2X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI2XL (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);



specify
if (B==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge S0 => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI2XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI4X1 (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(Y, YN);



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI4X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI4X2 (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(Y, YN);



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI4X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI4X4 (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(Y, YN);



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI4X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module MXI4XL (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(Y, YN);



specify
if (B==1'b0 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1 && D==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1 && D==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && D==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1)
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S1==1'b0)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S1==1'b1)
(S0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b1 && D==1'b1 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b0 && D==1'b1 && S0==1'b0)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1 && C==1'b1 && D==1'b0 && S0==1'b1)
(S1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // MXI4XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2BX1 (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2BX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2BX2 (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2BX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2BX4 (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2BX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2BXL (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2BXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2X1 (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2X2 (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2X4 (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND2XL (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND2XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BX1 (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (Y, Ax, B, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3BX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BX2 (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (Y, Ax, B, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3BX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BX4 (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (Y, Ax, B, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3BX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3BXL (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (Y, Ax, B, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3BXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3X1 (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3X2 (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3X4 (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND3XL (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND3XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BBX1 (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (Y, Ax, Bx, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BBX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BBX2 (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (Y, Ax, Bx, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BBX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BBX4 (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (Y, Ax, Bx, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BBX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BBXL (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nand (Y, Ax, Bx, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BBXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BX1 (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (Y, Ax, B, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BX2 (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (Y, Ax, B, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BX4 (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (Y, Ax, B, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4BXL (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (Y, Ax, B, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4BXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4X1 (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4X2 (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4X4 (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NAND4XL (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NAND4XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2BX1 (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2BX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2BX2 (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2BX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2BX4 (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2BX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2BXL (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor (Y, Ax, B);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2BXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2X1 (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2X2 (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2X4 (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR2XL (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR2XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BX1 (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nor (Y, Ax, B, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3BX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BX2 (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nor (Y, Ax, B, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3BX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BX4 (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nor (Y, Ax, B, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3BX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3BXL (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nor (Y, Ax, B, C);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3BXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3X1 (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3X2 (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3X4 (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR3XL (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR3XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BBX1 (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor (Y, Ax, Bx, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BBX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BBX2 (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor (Y, Ax, Bx, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BBX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BBX4 (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor (Y, Ax, Bx, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BBX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BBXL (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;

  not (Bx, BN);
  not (Ax, AN);
  nor (Y, Ax, Bx, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(BN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BBXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BX1 (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nor (Y, Ax, B, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BX2 (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nor (Y, Ax, B, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BX4 (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nor (Y, Ax, B, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4BXL (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nor (Y, Ax, B, C, D);


specify
(AN => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4BXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4X1 (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nor (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4X2 (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nor (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4X4 (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nor (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module NOR4XL (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nor (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // NOR4XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211X1 (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI211X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211X2 (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI211X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211X4 (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI211X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI211XL (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, C0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI211XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21X1 (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21X2 (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21X4 (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI21XL (Y, A0, A1, B0);
output Y;
input A0, A1, B0;



  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI21XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221X1 (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, C0, outB, outA);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI221X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221X2 (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, C0, outB, outA);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI221X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221X4 (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, C0, outB, outA);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI221X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI221XL (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, C0, outB, outA);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI221XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222X1 (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(Y, outA, outB, outC);


specify
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI222X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222X2 (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(Y, outA, outB, outC);


specify
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI222X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222X4 (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(Y, outA, outB, outC);


specify
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI222X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI222XL (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(Y, outA, outB, outC);


specify
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b0 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && C0==1'b1 && C1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b0 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && C0==1'b1 && C1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b0 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b0)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && B0==1'b1 && B1==1'b1)
(C1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI222XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22X1 (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22X2 (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22X4 (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI22XL (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;



  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI22XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB1X1 (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;



  nand I0 (outA, A0N, A1N);
  nand I1(Y, B0, outA);


specify
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2BB1X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB1X2 (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;



  nand I0 (outA, A0N, A1N);
  nand I1(Y, B0, outA);


specify
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2BB1X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB1X4 (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;



  nand I0 (outA, A0N, A1N);
  nand I1(Y, B0, outA);


specify
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2BB1X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB1XL (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;



  nand I0 (outA, A0N, A1N);
  nand I1(Y, B0, outA);


specify
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2BB1XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB2X1 (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;



  nand I0 (outA, A0N, A1N);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2BB2X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB2X2 (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;



  nand I0 (outA, A0N, A1N);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2BB2X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB2X4 (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;



  nand I0 (outA, A0N, A1N);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2BB2X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI2BB2XL (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;



  nand I0 (outA, A0N, A1N);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1N => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b0 && A1N==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0N==1'b1 && A1N==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI2BB2XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31X1 (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI31X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31X2 (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI31X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31X4 (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI31X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI31XL (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;



  or   I0(outA, A0, A1, A2);
  nand I1(Y, B0, outA);


specify
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI31XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI32X1 (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI32X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI32X2 (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI32X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI32X4 (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI32X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI32XL (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI32XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI33X1 (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1, B2);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI33X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI33X2 (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1, B2);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI33X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI33X4 (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1, B2);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI33X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OAI33XL (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;



  or   I0(outA, A0, A1, A2);
  or   I1(outB, B0, B1, B2);
  nand I2(Y, outA, outB);


specify
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b0 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b0 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b0)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B0==1'b1 && B1==1'b1 && B2==1'b1)
(A2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B0 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B1 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b0 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b0 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b0)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A0==1'b1 && A1==1'b1 && A2==1'b1)
(B2 => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OAI33XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2X1 (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2X2 (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2X4 (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR2XL (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR2XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3X1 (Y, A, B, C);
output Y;
input A, B, C;

  or (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3X2 (Y, A, B, C);
output Y;
input A, B, C;

  or (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3X4 (Y, A, B, C);
output Y;
input A, B, C;

  or (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR3XL (Y, A, B, C);
output Y;
input A, B, C;

  or (Y, A, B, C);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR3XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4X1 (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4X2 (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4X4 (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module OR4XL (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or (Y, A, B, C, D);


specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // OR4XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF1R1WX2 (RB, RW, RWN, WB, WW);
output RB;
input WB, WW, RW, RWN;
reg NOTIFIER;

   not II (wwn,WW);
   udp_tlatrf I0 (n0, WB, WW, wwn, NOTIFIER);
   notif1     I1 (RB, n0, n2);
   udp_outrf  I2 (n2, n0, RWN, RW);





wire ENABLE_RW_AND_NOT_RWN ;
assign ENABLE_RW_AND_NOT_RWN = (RW&!RWN) ? 1'b1:1'b0;

specify
(WB => RB) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WB==1'b0 && WW==1'b0)
( RW => RB ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WB==1'b1 && WW==1'b0)
( RW => RB ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WW==1'b1)
( RW => RB ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WB==1'b0 && WW==1'b0)
( RWN => RB ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WB==1'b1 && WW==1'b0)
( RWN => RB ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (WW==1'b1)
( RWN => RB ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge WW &&& (ENABLE_RW_AND_NOT_RWN == 1'b1), posedge WB, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WW &&& (ENABLE_RW_AND_NOT_RWN == 1'b1), negedge WB, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge WW &&& (ENABLE_RW_AND_NOT_RWN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge WW => (RB:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // RF1R1WX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RF2R1WX2 (R1B, R2B, R1W, R2W, WB, WW);
output R1B, R2B;
input WB, WW, R1W, R2W;
reg NOTIFIER;

   not        I0 (WWN, WW);
   not        I1 (R1WN, R1W);
   not        I2 (R2WN, R2W);
   udp_tlatrf I3 (n0, WB, WW, WWN, NOTIFIER);
   notif1     I4 (R1B, n0, n2);
   notif1     I5 (R2B, n0, n3);
   udp_outrf  I6 (n2, n0, R1WN, R1W);
   udp_outrf  I7 (n3, n0, R2WN, R2W);





wire ENABLE_R1W_OR_R2W ;
assign ENABLE_R1W_OR_R2W = (R1W | R2W) ? 1'b1:1'b0;

specify
if (R2W==1'b0)
(WB => R1B) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R2W==1'b1)
(WB => R1B) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R1W==1'b0)
(WB => R2B) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R1W==1'b1)
(WB => R2B) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R2W==1'b0 && WB==1'b0 && WW==1'b0)
( R1W => R1B ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R2W==1'b0 && WB==1'b1 && WW==1'b0)
( R1W => R1B ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R2W==1'b0 && WW==1'b1)
( R1W => R1B ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R2W==1'b1 && WB==1'b0 && WW==1'b0)
( R1W => R1B ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R2W==1'b1 && WB==1'b1 && WW==1'b0)
( R1W => R1B ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R2W==1'b1 && WW==1'b1)
( R1W => R1B ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R1W==1'b0 && WB==1'b0 && WW==1'b0)
( R2W => R2B ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R1W==1'b0 && WB==1'b1 && WW==1'b0)
( R2W => R2B ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R1W==1'b0 && WW==1'b1)
( R2W => R2B ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R1W==1'b1 && WB==1'b0 && WW==1'b0)
( R2W => R2B ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R1W==1'b1 && WB==1'b1 && WW==1'b0)
( R2W => R2B ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R1W==1'b1 && WW==1'b1)
( R2W => R2B ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge WW &&& (ENABLE_R1W_OR_R2W == 1'b1), posedge WB, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge WW &&& (ENABLE_R1W_OR_R2W == 1'b1), negedge WB, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge WW &&& (ENABLE_R1W_OR_R2W == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (R2W==1'b0)
(posedge WW => (R1B:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R2W==1'b1)
(posedge WW => (R1B:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R1W==1'b0)
(posedge WW => (R2B:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (R1W==1'b1)
(posedge WW => (R2B:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // RF2R1WX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RFRDX1 (BRB, RB);
output BRB;
input RB;
reg NOTIFIER;

   not(weak0,weak1) I0(RB, io_wire);
   not              I1(io_wire, RB);
   buf              I2(BRB, io_wire);






specify
(RB => BRB) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // RFRDX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RFRDX2 (BRB, RB);
output BRB;
input RB;
reg NOTIFIER;

   not(weak0,weak1) I0(RB, io_wire);
   not              I1(io_wire, RB);
   buf              I2(BRB, io_wire);






specify
(RB => BRB) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // RFRDX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RFRDX4 (BRB, RB);
output BRB;
input RB;
reg NOTIFIER;

   not(weak0,weak1) I0(RB, io_wire);
   not              I1(io_wire, RB);
   buf              I2(BRB, io_wire);






specify
(RB => BRB) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // RFRDX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RSLATNX1 (Q, QN, RN, SN);
output Q, QN;
input RN, SN;
reg NOTIFIER;
  not I4(R, RN);
  not I5(S, SN);
  udp_rslat  I0(q,  R, S, NOTIFIER);
  udp_rslatn I1(qn, R, S, NOTIFIER);
  not I2(QN, q);
  not I3(Q, qn);

wire ENABLE_SN ;
wire ENABLE_RN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge SN, posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (SN==1'b0)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (SN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // RSLATNX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RSLATNX2 (Q, QN, RN, SN);
output Q, QN;
input RN, SN;
reg NOTIFIER;
  not I4(R, RN);
  not I5(S, SN);
  udp_rslat  I0(q,  R, S, NOTIFIER);
  udp_rslatn I1(qn, R, S, NOTIFIER);
  not I2(QN, q);
  not I3(Q, qn);

wire ENABLE_SN ;
wire ENABLE_RN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge SN, posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (SN==1'b0)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (SN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // RSLATNX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RSLATNX4 (Q, QN, RN, SN);
output Q, QN;
input RN, SN;
reg NOTIFIER;
  not I4(R, RN);
  not I5(S, SN);
  udp_rslat  I0(q,  R, S, NOTIFIER);
  udp_rslatn I1(qn, R, S, NOTIFIER);
  not I2(QN, q);
  not I3(Q, qn);

wire ENABLE_SN ;
wire ENABLE_RN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge SN, posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (SN==1'b0)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (SN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // RSLATNX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RSLATNXL (Q, QN, RN, SN);
output Q, QN;
input RN, SN;
reg NOTIFIER;
  not I4(R, RN);
  not I5(S, SN);
  udp_rslat  I0(q,  R, S, NOTIFIER);
  udp_rslatn I1(qn, R, S, NOTIFIER);
  not I2(QN, q);
  not I3(Q, qn);

wire ENABLE_SN ;
wire ENABLE_RN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge SN, posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (SN==1'b0)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (SN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // RSLATNXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RSLATX1 (Q, QN, R, S);
output Q, QN;
input R, S;
reg NOTIFIER;
  udp_rslat  I0(q,  R, S, NOTIFIER);
  udp_rslatn I1(qn, R, S, NOTIFIER);
  buf I2(QN, qn);
  buf I3(Q, q);

wire ENABLE_NOT_S ;
wire ENABLE_NOT_R ;
assign ENABLE_NOT_S = (!S) ? 1'b1:1'b0;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;

specify
$width(posedge R &&& (ENABLE_NOT_S == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge S, negedge R, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R, negedge S, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge S &&& (ENABLE_NOT_R == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (S==1'b0)
(posedge R *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (S==1'b1)
(R => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (R==1'b0)
(posedge S *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (R==1'b1)
(S => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // RSLATX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RSLATX2 (Q, QN, R, S);
output Q, QN;
input R, S;
reg NOTIFIER;
  udp_rslat  I0(q,  R, S, NOTIFIER);
  udp_rslatn I1(qn, R, S, NOTIFIER);
  buf I2(QN, qn);
  buf I3(Q, q);

wire ENABLE_NOT_S ;
wire ENABLE_NOT_R ;
assign ENABLE_NOT_S = (!S) ? 1'b1:1'b0;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;

specify
$width(posedge R &&& (ENABLE_NOT_S == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge S, negedge R, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R, negedge S, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge S &&& (ENABLE_NOT_R == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (S==1'b0)
(posedge R *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (S==1'b1)
(R => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (R==1'b0)
(posedge S *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (R==1'b1)
(S => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // RSLATX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RSLATX4 (Q, QN, R, S);
output Q, QN;
input R, S;
reg NOTIFIER;
  udp_rslat  I0(q,  R, S, NOTIFIER);
  udp_rslatn I1(qn, R, S, NOTIFIER);
  buf I2(QN, qn);
  buf I3(Q, q);

wire ENABLE_NOT_S ;
wire ENABLE_NOT_R ;
assign ENABLE_NOT_S = (!S) ? 1'b1:1'b0;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;

specify
$width(posedge R &&& (ENABLE_NOT_S == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge S, negedge R, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R, negedge S, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge S &&& (ENABLE_NOT_R == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (S==1'b0)
(posedge R *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (S==1'b1)
(R => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (R==1'b0)
(posedge S *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (R==1'b1)
(S => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // RSLATX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module RSLATXL (Q, QN, R, S);
output Q, QN;
input R, S;
reg NOTIFIER;
  udp_rslat  I0(q,  R, S, NOTIFIER);
  udp_rslatn I1(qn, R, S, NOTIFIER);
  buf I2(QN, qn);
  buf I3(Q, q);

wire ENABLE_NOT_S ;
wire ENABLE_NOT_R ;
assign ENABLE_NOT_S = (!S) ? 1'b1:1'b0;
assign ENABLE_NOT_R = (!R) ? 1'b1:1'b0;

specify
$width(posedge R &&& (ENABLE_NOT_S == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge S, negedge R, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge R, negedge S, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge S &&& (ENABLE_NOT_R == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (S==1'b0)
(posedge R *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (S==1'b1)
(R => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
(posedge S *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(posedge R *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (R==1'b0)
(posedge S *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (R==1'b1)
(S => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // RSLATXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module SDFFHQX1 (Q, CK, D, SE, SI);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI = (D&!SI | !D&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFHQX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFHQX2 (Q, CK, D, SE, SI);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI = (D&!SI | !D&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFHQX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFHQX4 (Q, CK, D, SE, SI);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI = (D&!SI | !D&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFHQX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFHQXL (Q, CK, D, SE, SI);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI = (D&!SI | !D&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFHQXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNRX1 (Q, QN, CKN, D, RN, SE, SI);
output Q, QN;
input D, SI, SE, CKN, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI = (D&!SE | SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI = (D&RN&!SI | !D&RN&SI) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, negedge CKN &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // SDFFNRX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNRX2 (Q, QN, CKN, D, RN, SE, SI);
output Q, QN;
input D, SI, SE, CKN, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI = (D&!SE | SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI = (D&RN&!SI | !D&RN&SI) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, negedge CKN &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // SDFFNRX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNRX4 (Q, QN, CKN, D, RN, SE, SI);
output Q, QN;
input D, SI, SE, CKN, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI = (D&!SE | SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI = (D&RN&!SI | !D&RN&SI) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, negedge CKN &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // SDFFNRX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNRXL (Q, QN, CKN, D, RN, SE, SI);
output Q, QN;
input D, SI, SE, CKN, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI = (D&!SE | SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI = (D&RN&!SI | !D&RN&SI) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, negedge CKN &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // SDFFNRXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSRX1 (Q, QN, CKN, D, RN, SE, SI, SN);
output Q, QN;
input D, SI, SE, CKN, SN, RN;
reg NOTIFIER;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN = (D&!SE&SN | SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN = (D&RN&!SI&SN | !D&RN&SI&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI = (!D&RN&!SE | RN&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNSRX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSRX2 (Q, QN, CKN, D, RN, SE, SI, SN);
output Q, QN;
input D, SI, SE, CKN, SN, RN;
reg NOTIFIER;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN = (D&!SE&SN | SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN = (D&RN&!SI&SN | !D&RN&SI&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI = (!D&RN&!SE | RN&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNSRX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSRX4 (Q, QN, CKN, D, RN, SE, SI, SN);
output Q, QN;
input D, SI, SE, CKN, SN, RN;
reg NOTIFIER;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN = (D&!SE&SN | SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN = (D&RN&!SI&SN | !D&RN&SI&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI = (!D&RN&!SE | RN&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNSRX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSRXL (Q, QN, CKN, D, RN, SE, SI, SN);
output Q, QN;
input D, SI, SE, CKN, SN, RN;
reg NOTIFIER;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN = (D&!SE&SN | SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN = (D&RN&!SI&SN | !D&RN&SI&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI = (!D&RN&!SE | RN&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, negedge CKN &&& (ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNSRXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSX1 (Q, QN, CKN, D, SE, SI, SN);
output Q, QN;
input D, SI, SE, CKN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN ;
wire ENABLE_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN = (D&!SI&SN | !D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI = (!D&!SE | SE&!SI) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNSX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSX2 (Q, QN, CKN, D, SE, SI, SN);
output Q, QN;
input D, SI, SE, CKN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN ;
wire ENABLE_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN = (D&!SI&SN | !D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI = (!D&!SE | SE&!SI) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNSX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSX4 (Q, QN, CKN, D, SE, SI, SN);
output Q, QN;
input D, SI, SE, CKN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN ;
wire ENABLE_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN = (D&!SI&SN | !D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI = (!D&!SE | SE&!SI) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNSX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNSXL (Q, QN, CKN, D, SE, SI, SN);
output Q, QN;
input D, SI, SE, CKN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN ;
wire ENABLE_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN = (D&!SI&SN | !D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI = (!D&!SE | SE&!SI) ? 1'b1:1'b0;

specify
$width(posedge CKN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CKN==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFNSXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNX1 (Q, QN, CKN, D, SE, SI);
output Q, QN;
input D, SI, SE, CKN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI = (D&!SI | !D&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CKN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFNX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNX2 (Q, QN, CKN, D, SE, SI);
output Q, QN;
input D, SI, SE, CKN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI = (D&!SI | !D&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CKN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFNX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNX4 (Q, QN, CKN, D, SE, SI);
output Q, QN;
input D, SI, SE, CKN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI = (D&!SI | !D&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CKN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFNX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFNXL (Q, QN, CKN, D, SE, SI);
output Q, QN;
input D, SI, SE, CKN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, CKN);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI = (D&!SI | !D&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CKN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CKN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(negedge CKN => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFNXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRHQX1 (Q, CK, D, RN, SE, SI);
output Q;
input D, SI, SE, CK, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI = (D&!SE | SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI = (D&RN&!SI | !D&RN&SI) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFRHQX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRHQX2 (Q, CK, D, RN, SE, SI);
output Q;
input D, SI, SE, CK, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI = (D&!SE | SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI = (D&RN&!SI | !D&RN&SI) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFRHQX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRHQX4 (Q, CK, D, RN, SE, SI);
output Q;
input D, SI, SE, CK, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI = (D&!SE | SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI = (D&RN&!SI | !D&RN&SI) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFRHQX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRHQXL (Q, CK, D, RN, SE, SI);
output Q;
input D, SI, SE, CK, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI = (D&!SE | SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI = (D&RN&!SI | !D&RN&SI) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFRHQXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRX1 (Q, QN, CK, D, RN, SE, SI);
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI = (D&!SE | SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI = (D&RN&!SI | !D&RN&SI) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // SDFFRX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRX2 (Q, QN, CK, D, RN, SE, SI);
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI = (D&!SE | SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI = (D&RN&!SI | !D&RN&SI) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // SDFFRX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRX4 (Q, QN, CK, D, RN, SE, SI);
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI = (D&!SE | SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI = (D&RN&!SI | !D&RN&SI) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // SDFFRX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFRXL (Q, QN, CK, D, RN, SE, SI);
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI ;
wire ENABLE_RN_AND_SE ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI = (D&!SE | SE&SI) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI = (D&RN&!SI | !D&RN&SI) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE = (RN&SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // SDFFRXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSHQX1 (Q, CK, D, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN ;
wire ENABLE_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN = (D&!SI&SN | !D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI = (!D&!SE | SE&!SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // SDFFSHQX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSHQX2 (Q, CK, D, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN ;
wire ENABLE_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN = (D&!SI&SN | !D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI = (!D&!SE | SE&!SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // SDFFSHQX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSHQX4 (Q, CK, D, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN ;
wire ENABLE_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN = (D&!SI&SN | !D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI = (!D&!SE | SE&!SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // SDFFSHQX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSHQXL (Q, CK, D, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN ;
wire ENABLE_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN = (D&!SI&SN | !D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI = (!D&!SE | SE&!SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // SDFFSHQXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRHQX1 (Q, CK, D, RN, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN = (D&!SE&SN | SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN = (D&RN&!SI&SN | !D&RN&SI&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI = (!D&RN&!SE | RN&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // SDFFSRHQX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRHQX2 (Q, CK, D, RN, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN = (D&!SE&SN | SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN = (D&RN&!SI&SN | !D&RN&SI&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI = (!D&RN&!SE | RN&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // SDFFSRHQX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRHQX4 (Q, CK, D, RN, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN = (D&!SE&SN | SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN = (D&RN&!SI&SN | !D&RN&SI&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI = (!D&RN&!SE | RN&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // SDFFSRHQX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRHQXL (Q, CK, D, RN, SE, SI, SN);
output Q;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN = (D&!SE&SN | SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN = (D&RN&!SI&SN | !D&RN&SI&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI = (!D&RN&!SE | RN&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // SDFFSRHQXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRX1 (Q, QN, CK, D, RN, SE, SI, SN);
output Q, QN;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN = (D&!SE&SN | SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN = (D&RN&!SI&SN | !D&RN&SI&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI = (!D&RN&!SE | RN&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSRX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRX2 (Q, QN, CK, D, RN, SE, SI, SN);
output Q, QN;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN = (D&!SE&SN | SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN = (D&RN&!SI&SN | !D&RN&SI&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI = (!D&RN&!SE | RN&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSRX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRX4 (Q, QN, CK, D, RN, SE, SI, SN);
output Q, QN;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN = (D&!SE&SN | SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN = (D&RN&!SI&SN | !D&RN&SI&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI = (!D&RN&!SE | RN&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSRX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSRXL (Q, QN, CK, D, RN, SE, SI, SN);
output Q, QN;
input D, SI, SE, CK, SN, RN;
reg NOTIFIER;
  buf   XX0 (xRN, RN);
  buf   XX1 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_RN_AND_SN ;
wire ENABLE_RN_AND_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN ;
wire ENABLE_SN ;
wire ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN ;
wire ENABLE_RN_AND_SE_AND_SN ;
wire ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI ;
wire ENABLE_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE_AND_SN = (RN&!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN = (D&!SE&SN | SE&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN = (D&RN&!SI&SN | !D&RN&SI&SN) ? 1'b1:1'b0;
assign ENABLE_RN_AND_SE_AND_SN = (RN&SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI = (!D&RN&!SE | RN&SE&!SI) ? 1'b1:1'b0;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge RN, posedge CK &&& (ENABLE_D_AND_NOT_SE_AND_SN_OR_SE_AND_SI_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_AND_SN_OR_NOT_D_AND_RN_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_RN_AND_NOT_SE_OR_RN_AND_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN, posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSRXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSX1 (Q, QN, CK, D, SE, SI, SN);
output Q, QN;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN ;
wire ENABLE_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN = (D&!SI&SN | !D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI = (!D&!SE | SE&!SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSX2 (Q, QN, CK, D, SE, SI, SN);
output Q, QN;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN ;
wire ENABLE_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN = (D&!SI&SN | !D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI = (!D&!SE | SE&!SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSX4 (Q, QN, CK, D, SE, SI, SN);
output Q, QN;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN ;
wire ENABLE_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN = (D&!SI&SN | !D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI = (!D&!SE | SE&!SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFSXL (Q, QN, CK, D, SE, SI, SN);
output Q, QN;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_SN ;
wire ENABLE_NOT_SE_AND_SN ;
wire ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN ;
wire ENABLE_SE_AND_SN ;
wire ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_SE_AND_SN = (!SE&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN = (D&!SI&SN | !D&SI&SN) ? 1'b1:1'b0;
assign ENABLE_SE_AND_SN = (SE&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI = (!D&!SE | SE&!SI) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_AND_SN_OR_NOT_D_AND_SI_AND_SN == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE_AND_SN == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$recrem(posedge SN, posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b0 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b0 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b0 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (CK==1'b1 && D==1'b1 && SE==1'b1 && SI==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // SDFFSXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFTRX1 (Q, QN, CK, D, RN, SE, SI);
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
   udp_sedfft I0 (n0, D, CK, xRN, SI, SE, 1'b1, NOTIFIER);
   buf        I1 (Q, n0);
   not        I2 (QN, n0);

wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_RN_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE = (D&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_RN_AND_SI = (D&RN&!SI | !D&SI | !RN&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFTRX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFTRX2 (Q, QN, CK, D, RN, SE, SI);
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
   udp_sedfft I0 (n0, D, CK, xRN, SI, SE, 1'b1, NOTIFIER);
   buf        I1 (Q, n0);
   not        I2 (QN, n0);

wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_RN_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE = (D&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_RN_AND_SI = (D&RN&!SI | !D&SI | !RN&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFTRX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFTRX4 (Q, QN, CK, D, RN, SE, SI);
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
   udp_sedfft I0 (n0, D, CK, xRN, SI, SE, 1'b1, NOTIFIER);
   buf        I1 (Q, n0);
   not        I2 (QN, n0);

wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_RN_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE = (D&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_RN_AND_SI = (D&RN&!SI | !D&SI | !RN&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFTRX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFTRXL (Q, QN, CK, D, RN, SE, SI);
output Q, QN;
input D, SI, SE, CK, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  buf   XX0 (xRN, RN);
   udp_sedfft I0 (n0, D, CK, xRN, SI, SE, 1'b1, NOTIFIER);
   buf        I1 (Q, n0);
   not        I2 (QN, n0);

wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_RN_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE = (D&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_RN_AND_SI = (D&RN&!SI | !D&SI | !RN&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && RN==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFTRXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFX1 (Q, QN, CK, D, SE, SI);
output Q, QN;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI = (D&!SI | !D&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFX1
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFX2 (Q, QN, CK, D, SE, SI);
output Q, QN;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI = (D&!SI | !D&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFX2
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFX4 (Q, QN, CK, D, SE, SI);
output Q, QN;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI = (D&!SI | !D&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFX4
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SDFFXL (Q, QN, CK, D, SE, SI);
output Q, QN;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
  udp_mux2 I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  not     I72 (QN, n0);

wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI = (D&!SI | !D&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SDFFXL
`endcelldefine
	

`timescale 1ns/1ps
`celldefine
module SEDFFHQX1 (Q, CK, D, E, SE, SI);
output Q;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR I0 (n0, D, CK, xRN, SI, SE, E, 1'b1, 1'b0, NOTIFIER);
   buf       I1 (Q, n0);

wire ENABLE_E_OR_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E ;
wire ENABLE_SE ;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E = (D&!SI | !D&SI | !E) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFHQX1
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFHQX2 (Q, CK, D, E, SE, SI);
output Q;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR I0 (n0, D, CK, xRN, SI, SE, E, 1'b1, 1'b0, NOTIFIER);
   buf       I1 (Q, n0);

wire ENABLE_E_OR_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E ;
wire ENABLE_SE ;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E = (D&!SI | !D&SI | !E) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFHQX2
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFHQX4 (Q, CK, D, E, SE, SI);
output Q;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR I0 (n0, D, CK, xRN, SI, SE, E, 1'b1, 1'b0, NOTIFIER);
   buf       I1 (Q, n0);

wire ENABLE_E_OR_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E ;
wire ENABLE_SE ;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E = (D&!SI | !D&SI | !E) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFHQX4
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFHQXL (Q, CK, D, E, SE, SI);
output Q;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR I0 (n0, D, CK, xRN, SI, SE, E, 1'b1, 1'b0, NOTIFIER);
   buf       I1 (Q, n0);

wire ENABLE_E_OR_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E ;
wire ENABLE_SE ;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E = (D&!SI | !D&SI | !E) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFHQXL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFTRX1 (Q, QN, CK, D, E, RN, SE, SI);
output Q, QN;
input D, CK, E, SE, SI, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

   udp_sedfft I0 (n0, D, CK, xRN, SI, SE, E, NOTIFIER);
   buf        I1 (Q, n0);
   not        I2 (QN, n0);

wire ENABLE_E_OR_NOT_RN_OR_SE ;
wire ENABLE_E_AND_RN_AND_NOT_SE ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE_OR_NOT_E_AND_NOT_SE ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E_AND_RN_OR_NOT_RN_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_E_OR_NOT_RN_OR_SE = (E | !RN | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_RN_AND_NOT_SE = (E&RN&!SE) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_OR_NOT_E_AND_NOT_SE = (D&!SE | !E&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E_AND_RN_OR_NOT_RN_AND_SI = (D&RN&!SI | !D&SI | !E&RN | !RN&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_NOT_RN_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_NOT_RN_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_NOT_E_AND_NOT_SE == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_NOT_E_AND_NOT_SE == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E_AND_RN_OR_NOT_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E_AND_RN_OR_NOT_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFTRX1
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFTRX2 (Q, QN, CK, D, E, RN, SE, SI);
output Q, QN;
input D, CK, E, SE, SI, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

   udp_sedfft I0 (n0, D, CK, xRN, SI, SE, E, NOTIFIER);
   buf        I1 (Q, n0);
   not        I2 (QN, n0);

wire ENABLE_E_OR_NOT_RN_OR_SE ;
wire ENABLE_E_AND_RN_AND_NOT_SE ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE_OR_NOT_E_AND_NOT_SE ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E_AND_RN_OR_NOT_RN_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_E_OR_NOT_RN_OR_SE = (E | !RN | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_RN_AND_NOT_SE = (E&RN&!SE) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_OR_NOT_E_AND_NOT_SE = (D&!SE | !E&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E_AND_RN_OR_NOT_RN_AND_SI = (D&RN&!SI | !D&SI | !E&RN | !RN&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_NOT_RN_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_NOT_RN_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_NOT_E_AND_NOT_SE == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_NOT_E_AND_NOT_SE == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E_AND_RN_OR_NOT_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E_AND_RN_OR_NOT_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFTRX2
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFTRX4 (Q, QN, CK, D, E, RN, SE, SI);
output Q, QN;
input D, CK, E, SE, SI, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

   udp_sedfft I0 (n0, D, CK, xRN, SI, SE, E, NOTIFIER);
   buf        I1 (Q, n0);
   not        I2 (QN, n0);

wire ENABLE_E_OR_NOT_RN_OR_SE ;
wire ENABLE_E_AND_RN_AND_NOT_SE ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE_OR_NOT_E_AND_NOT_SE ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E_AND_RN_OR_NOT_RN_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_E_OR_NOT_RN_OR_SE = (E | !RN | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_RN_AND_NOT_SE = (E&RN&!SE) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_OR_NOT_E_AND_NOT_SE = (D&!SE | !E&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E_AND_RN_OR_NOT_RN_AND_SI = (D&RN&!SI | !D&SI | !E&RN | !RN&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_NOT_RN_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_NOT_RN_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_NOT_E_AND_NOT_SE == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_NOT_E_AND_NOT_SE == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E_AND_RN_OR_NOT_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E_AND_RN_OR_NOT_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFTRX4
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFTRXL (Q, QN, CK, D, E, RN, SE, SI);
output Q, QN;
input D, CK, E, SE, SI, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;
  buf   XX1 (xRN, RN);

   udp_sedfft I0 (n0, D, CK, xRN, SI, SE, E, NOTIFIER);
   buf        I1 (Q, n0);
   not        I2 (QN, n0);

wire ENABLE_E_OR_NOT_RN_OR_SE ;
wire ENABLE_E_AND_RN_AND_NOT_SE ;
wire ENABLE_RN_AND_NOT_SE ;
wire ENABLE_D_AND_NOT_SE_OR_NOT_E_AND_NOT_SE ;
wire ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E_AND_RN_OR_NOT_RN_AND_SI ;
wire ENABLE_SE ;
assign ENABLE_E_OR_NOT_RN_OR_SE = (E | !RN | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_RN_AND_NOT_SE = (E&RN&!SE) ? 1'b1:1'b0;
assign ENABLE_RN_AND_NOT_SE = (RN&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SE_OR_NOT_E_AND_NOT_SE = (D&!SE | !E&!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E_AND_RN_OR_NOT_RN_AND_SI = (D&RN&!SI | !D&SI | !E&RN | !RN&SI) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_NOT_RN_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_NOT_RN_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_RN_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_RN_AND_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_NOT_E_AND_NOT_SE == 1'b1), posedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_NOT_E_AND_NOT_SE == 1'b1), negedge RN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E_AND_RN_OR_NOT_RN_AND_SI == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_RN_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E_AND_RN_OR_NOT_RN_AND_SI == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && RN==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b0 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b0 && RN==1'b0 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && RN==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && RN==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFTRXL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFX1 (Q, QN, CK, D, E, SE, SI);
output Q, QN;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR I0 (n0, D, CK, xRN, SI, SE, E, 1'b1, 1'b0, NOTIFIER); 
  buf     I1 (Q, n0);  
  not     I2 (QN, n0);

wire ENABLE_E_OR_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E ;
wire ENABLE_SE ;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E = (D&!SI | !D&SI | !E) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFX1
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFX2 (Q, QN, CK, D, E, SE, SI);
output Q, QN;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR I0 (n0, D, CK, xRN, SI, SE, E, 1'b1, 1'b0, NOTIFIER); 
  buf     I1 (Q, n0);  
  not     I2 (QN, n0);

wire ENABLE_E_OR_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E ;
wire ENABLE_SE ;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E = (D&!SI | !D&SI | !E) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFX2
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFX4 (Q, QN, CK, D, E, SE, SI);
output Q, QN;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR I0 (n0, D, CK, xRN, SI, SE, E, 1'b1, 1'b0, NOTIFIER); 
  buf     I1 (Q, n0);  
  not     I2 (QN, n0);

wire ENABLE_E_OR_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E ;
wire ENABLE_SE ;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E = (D&!SI | !D&SI | !E) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFX4
`endcelldefine


`timescale 1ns/1ps
`celldefine
module SEDFFXL (Q, QN, CK, D, E, SE, SI);
output Q, QN;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff_PWR I0 (n0, D, CK, xRN, SI, SE, E, 1'b1, 1'b0, NOTIFIER); 
  buf     I1 (Q, n0);  
  not     I2 (QN, n0);

wire ENABLE_E_OR_SE ;
wire ENABLE_E_AND_NOT_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E ;
wire ENABLE_SE ;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_E_AND_NOT_SE = (E&!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E = (D&!SI | !D&SI | !E) ? 1'b1:1'b0;
assign ENABLE_SE = (SE) ? 1'b1:1'b0;

specify
$width(posedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SI_OR_NOT_D_AND_SI_OR_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), posedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_SE == 1'b1), negedge SI, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b0 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && E==1'b1 && SI==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b1 || D==1'b0 && E==1'b1 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b0 && SI==1'b1 || D==1'b1 && E==1'b0 && SE==1'b1 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && E==1'b1 && SE==1'b1)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0 && SI==1'b0)
(posedge CK => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // SEDFFXL
`endcelldefine


`timescale 1ns/1ps
`celldefine
module TBUFIX1 (Y, A, OE);
output Y;
input A, OE;

  notif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFIX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFIX12 (Y, A, OE);
output Y;
input A, OE;

  notif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFIX12
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFIX16 (Y, A, OE);
output Y;
input A, OE;

  notif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFIX16
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFIX2 (Y, A, OE);
output Y;
input A, OE;

  notif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFIX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFIX20 (Y, A, OE);
output Y;
input A, OE;

  notif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFIX20
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFIX3 (Y, A, OE);
output Y;
input A, OE;

  notif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFIX3
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFIX4 (Y, A, OE);
output Y;
input A, OE;

  notif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFIX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFIX8 (Y, A, OE);
output Y;
input A, OE;

  notif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFIX8
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFIXL (Y, A, OE);
output Y;
input A, OE;

  notif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFIXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFX1 (Y, A, OE);
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFX12 (Y, A, OE);
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFX12
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFX16 (Y, A, OE);
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFX16
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFX2 (Y, A, OE);
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFX20 (Y, A, OE);
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFX20
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFX3 (Y, A, OE);
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFX3
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFX4 (Y, A, OE);
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFX8 (Y, A, OE);
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFX8
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TBUFXL (Y, A, OE);
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);



specify
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
( OE => Y ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TBUFXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TIEHI (Y);
output Y;

  buf I0(Y, 1'b1);


specify

endspecify
endmodule // TIEHI
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TIELO (Y);
output Y;

  buf I0(Y, 1'b0);


specify

endspecify
endmodule // TIELO
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATCOX1 (ECKN, CKN, E);
output ECKN;
input  E, CKN;
reg NOTIFIER;

supply1 R, S;

  not      I0 (nclk,CKN);
  udp_tlat_PWR I1 (n0, E, nclk, R, S, 1'b1, 1'b0, NOTIFIER);
  not      I2 (nn0,n0);
  or       I3 (ECKN, nn0, CKN);


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CKN => ECKN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(posedge CKN => (ECKN:1'bx)) = (`ARM_PROP_DELAY,`ARM_INVALID_DELAY);
$width(posedge CKN &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(posedge CKN &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATCOX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATCOX2 (ECKN, CKN, E);
output ECKN;
input  E, CKN;
reg NOTIFIER;

supply1 R, S;

  not      I0 (nclk,CKN);
  udp_tlat_PWR I1 (n0, E, nclk, R, S, 1'b1, 1'b0, NOTIFIER);
  not      I2 (nn0,n0);
  or       I3 (ECKN, nn0, CKN);


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CKN => ECKN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(posedge CKN => (ECKN:1'bx)) = (`ARM_PROP_DELAY,`ARM_INVALID_DELAY);
$width(posedge CKN &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(posedge CKN &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATCOX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATCOX3 (ECKN, CKN, E);
output ECKN;
input  E, CKN;
reg NOTIFIER;

supply1 R, S;

  not      I0 (nclk,CKN);
  udp_tlat_PWR I1 (n0, E, nclk, R, S, 1'b1, 1'b0, NOTIFIER);
  not      I2 (nn0,n0);
  or       I3 (ECKN, nn0, CKN);


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CKN => ECKN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(posedge CKN => (ECKN:1'bx)) = (`ARM_PROP_DELAY,`ARM_INVALID_DELAY);
$width(posedge CKN &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(posedge CKN &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATCOX3
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATCOX4 (ECKN, CKN, E);
output ECKN;
input  E, CKN;
reg NOTIFIER;

supply1 R, S;

  not      I0 (nclk,CKN);
  udp_tlat_PWR I1 (n0, E, nclk, R, S, 1'b1, 1'b0, NOTIFIER);
  not      I2 (nn0,n0);
  or       I3 (ECKN, nn0, CKN);


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CKN => ECKN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(posedge CKN => (ECKN:1'bx)) = (`ARM_PROP_DELAY,`ARM_INVALID_DELAY);
$width(posedge CKN &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(posedge CKN &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATCOX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNCAX1 (ECK, CK, E);
output ECK;
input  E, CK;
reg NOTIFIER;

supply1 R, S;

  udp_tlat_PWR I0 (n0, E, CK, R, S, 1'b1, 1'b0, NOTIFIER);
  and      I1 (ECK, n0, CK);


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(negedge CK => (ECK:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATNCAX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNCAX2 (ECK, CK, E);
output ECK;
input  E, CK;
reg NOTIFIER;

supply1 R, S;

  udp_tlat_PWR I0 (n0, E, CK, R, S, 1'b1, 1'b0, NOTIFIER);
  and      I1 (ECK, n0, CK);


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(negedge CK => (ECK:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATNCAX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNCAX3 (ECK, CK, E);
output ECK;
input  E, CK;
reg NOTIFIER;

supply1 R, S;

  udp_tlat_PWR I0 (n0, E, CK, R, S, 1'b1, 1'b0, NOTIFIER);
  and      I1 (ECK, n0, CK);


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(negedge CK => (ECK:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATNCAX3
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNCAX4 (ECK, CK, E);
output ECK;
input  E, CK;
reg NOTIFIER;

supply1 R, S;

  udp_tlat_PWR I0 (n0, E, CK, R, S, 1'b1, 1'b0, NOTIFIER);
  and      I1 (ECK, n0, CK);


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(negedge CK => (ECK:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATNCAX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNCAX6 (ECK, CK, E);
output ECK;
input  E, CK;
reg NOTIFIER;

supply1 R, S;

  udp_tlat_PWR I0 (n0, E, CK, R, S, 1'b1, 1'b0, NOTIFIER);
  and      I1 (ECK, n0, CK);


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(negedge CK => (ECK:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATNCAX6
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNCAX8 (ECK, CK, E);
output ECK;
input  E, CK;
reg NOTIFIER;

supply1 R, S;

  udp_tlat_PWR I0 (n0, E, CK, R, S, 1'b1, 1'b0, NOTIFIER);
  and      I1 (ECK, n0, CK);


wire ENABLE_NOT_E ;
wire ENABLE_E ;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
assign ENABLE_E = (E) ? 1'b1:1'b0;

specify
if (E==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0)
(negedge CK => (ECK:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK, posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK, negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATNCAX8
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNRX1 (Q, QN, D, GN, RN);
output  Q, QN;
input  D, GN, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, GN);

wire ENABLE_RN ;
wire ENABLE_D ;
wire ENABLE_GN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_GN = (GN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge RN, posedge GN &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_GN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // TLATNRX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNRX2 (Q, QN, D, GN, RN);
output  Q, QN;
input  D, GN, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, GN);

wire ENABLE_RN ;
wire ENABLE_D ;
wire ENABLE_GN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_GN = (GN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge RN, posedge GN &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_GN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // TLATNRX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNRX4 (Q, QN, D, GN, RN);
output  Q, QN;
input  D, GN, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, GN);

wire ENABLE_RN ;
wire ENABLE_D ;
wire ENABLE_GN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_GN = (GN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge RN, posedge GN &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_GN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // TLATNRX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNRXL (Q, QN, D, GN, RN);
output  Q, QN;
input  D, GN, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, GN);

wire ENABLE_RN ;
wire ENABLE_D ;
wire ENABLE_GN ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_GN = (GN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge RN, posedge GN &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_GN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);

endspecify
endmodule // TLATNRXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNSRX1 (Q, QN, D, GN, RN, SN);
output  Q, QN;
input  D, GN, RN, SN;
reg NOTIFIER;

buf       XX0 (xSN, SN);
buf       XX1 (xRN, RN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_GN_AND_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_GN ;
wire ENABLE_GN_AND_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_GN_AND_SN = (GN&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_GN = (GN) ? 1'b1:1'b0;
assign ENABLE_GN_AND_RN = (GN&RN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge RN, posedge GN &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_GN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge GN &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN &&& (ENABLE_GN == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_GN_AND_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && GN==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATNSRX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNSRX2 (Q, QN, D, GN, RN, SN);
output  Q, QN;
input  D, GN, RN, SN;
reg NOTIFIER;

buf       XX0 (xSN, SN);
buf       XX1 (xRN, RN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_GN_AND_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_GN ;
wire ENABLE_GN_AND_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_GN_AND_SN = (GN&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_GN = (GN) ? 1'b1:1'b0;
assign ENABLE_GN_AND_RN = (GN&RN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge RN, posedge GN &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_GN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge GN &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN &&& (ENABLE_GN == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_GN_AND_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && GN==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATNSRX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNSRX4 (Q, QN, D, GN, RN, SN);
output  Q, QN;
input  D, GN, RN, SN;
reg NOTIFIER;

buf       XX0 (xSN, SN);
buf       XX1 (xRN, RN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_GN_AND_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_GN ;
wire ENABLE_GN_AND_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_GN_AND_SN = (GN&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_GN = (GN) ? 1'b1:1'b0;
assign ENABLE_GN_AND_RN = (GN&RN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge RN, posedge GN &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_GN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge GN &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN &&& (ENABLE_GN == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_GN_AND_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && GN==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATNSRX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNSRXL (Q, QN, D, GN, RN, SN);
output  Q, QN;
input  D, GN, RN, SN;
reg NOTIFIER;

buf       XX0 (xSN, SN);
buf       XX1 (xRN, RN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_GN_AND_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_GN ;
wire ENABLE_GN_AND_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_GN_AND_SN = (GN&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_GN = (GN) ? 1'b1:1'b0;
assign ENABLE_GN_AND_RN = (GN&RN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge RN, posedge GN &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_GN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge GN &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN &&& (ENABLE_GN == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_GN_AND_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && GN==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && GN==1'b0)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0 && RN==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATNSRXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNSX1 (Q, QN, D, GN, SN);
output  Q, QN;
input  D, GN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, GN);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_GN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_GN = (GN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_GN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATNSX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNSX2 (Q, QN, D, GN, SN);
output  Q, QN;
input  D, GN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, GN);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_GN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_GN = (GN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_GN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATNSX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNSX4 (Q, QN, D, GN, SN);
output  Q, QN;
input  D, GN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, GN);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_GN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_GN = (GN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_GN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATNSX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNSXL (Q, QN, D, GN, SN);
output  Q, QN;
input  D, GN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, GN);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_GN ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_GN = (GN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, posedge GN &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_GN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && GN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATNSXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNTSCAX1 (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR I1 (n0, n1, CK, R, S, 1'b1, 1'b0, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATNTSCAX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNTSCAX2 (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR I1 (n0, n1, CK, R, S, 1'b1, 1'b0, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATNTSCAX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNTSCAX3 (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR I1 (n0, n1, CK, R, S, 1'b1, 1'b0, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATNTSCAX3
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNTSCAX4 (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR I1 (n0, n1, CK, R, S, 1'b1, 1'b0, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATNTSCAX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNTSCAX6 (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR I1 (n0, n1, CK, R, S, 1'b1, 1'b0, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATNTSCAX6
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNTSCAX8 (ECK, CK, E, SE);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat_PWR I1 (n0, n1, CK, R, S, 1'b1, 1'b0, NOTIFIER);
  and      I2 (ECK, n0, CK);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CK => ECK) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(negedge CK => (ECK:1'bx)) = (`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
$width(negedge CK &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(negedge CK &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge CK &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATNTSCAX8
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNX1 (Q, QN, D, GN);
output  Q, QN;
input  D, GN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);


specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TLATNX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNX2 (Q, QN, D, GN);
output  Q, QN;
input  D, GN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);


specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TLATNX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNX4 (Q, QN, D, GN);
output  Q, QN;
input  D, GN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);


specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TLATNX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATNXL (Q, QN, D, GN);
output  Q, QN;
input  D, GN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);


specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(posedge GN, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(posedge GN, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge GN,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(negedge GN => (Q:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge GN => (QN:1'bx))=(`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TLATNXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATRX1 (Q, QN, D, G, RN);
output  Q, QN;
input  D, G, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_RN ;
wire ENABLE_D ;
wire ENABLE_NOT_G ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_G = (!G) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge RN, negedge G &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_NOT_G == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b1)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATRX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATRX2 (Q, QN, D, G, RN);
output  Q, QN;
input  D, G, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_RN ;
wire ENABLE_D ;
wire ENABLE_NOT_G ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_G = (!G) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge RN, negedge G &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_NOT_G == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b1)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATRX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATRX4 (Q, QN, D, G, RN);
output  Q, QN;
input  D, G, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_RN ;
wire ENABLE_D ;
wire ENABLE_NOT_G ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_G = (!G) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge RN, negedge G &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_NOT_G == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b1)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATRX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATRXL (Q, QN, D, G, RN);
output  Q, QN;
input  D, G, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_RN ;
wire ENABLE_D ;
wire ENABLE_NOT_G ;
assign ENABLE_RN = (RN) ? 1'b1:1'b0;
assign ENABLE_D = (D) ? 1'b1:1'b0;
assign ENABLE_NOT_G = (!G) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_RN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_RN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge RN, negedge G &&& (ENABLE_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_NOT_G == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b1)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATRXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATSRX1 (Q, QN, D, G, RN, SN);
output  Q, QN;
input  D, G, SN, RN;
reg NOTIFIER;

buf       XX0 (xSN, SN);
buf       XX1 (xRN, RN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_G_AND_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_NOT_G ;
wire ENABLE_NOT_G_AND_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_G_AND_SN = (!G&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_NOT_G = (!G) ? 1'b1:1'b0;
assign ENABLE_NOT_G_AND_RN = (!G&RN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge RN, negedge G &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_NOT_G_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, negedge G &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN &&& (ENABLE_NOT_G == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_G_AND_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b1)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATSRX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATSRX2 (Q, QN, D, G, RN, SN);
output  Q, QN;
input  D, G, SN, RN;
reg NOTIFIER;

buf       XX0 (xSN, SN);
buf       XX1 (xRN, RN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_G_AND_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_NOT_G ;
wire ENABLE_NOT_G_AND_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_G_AND_SN = (!G&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_NOT_G = (!G) ? 1'b1:1'b0;
assign ENABLE_NOT_G_AND_RN = (!G&RN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge RN, negedge G &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_NOT_G_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, negedge G &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN &&& (ENABLE_NOT_G == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_G_AND_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b1)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATSRX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATSRX4 (Q, QN, D, G, RN, SN);
output  Q, QN;
input  D, G, SN, RN;
reg NOTIFIER;

buf       XX0 (xSN, SN);
buf       XX1 (xRN, RN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_G_AND_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_NOT_G ;
wire ENABLE_NOT_G_AND_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_G_AND_SN = (!G&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_NOT_G = (!G) ? 1'b1:1'b0;
assign ENABLE_NOT_G_AND_RN = (!G&RN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge RN, negedge G &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_NOT_G_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, negedge G &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN &&& (ENABLE_NOT_G == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_G_AND_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b1)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATSRX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATSRXL (Q, QN, D, G, RN, SN);
output  Q, QN;
input  D, G, SN, RN;
reg NOTIFIER;

buf       XX0 (xSN, SN);
buf       XX1 (xRN, RN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_RN_AND_SN ;
wire ENABLE_D_AND_SN ;
wire ENABLE_NOT_G_AND_SN ;
wire ENABLE_NOT_D_AND_RN ;
wire ENABLE_NOT_G ;
wire ENABLE_NOT_G_AND_RN ;
assign ENABLE_RN_AND_SN = (RN&SN) ? 1'b1:1'b0;
assign ENABLE_D_AND_SN = (D&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_G_AND_SN = (!G&SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D_AND_RN = (!D&RN) ? 1'b1:1'b0;
assign ENABLE_NOT_G = (!G) ? 1'b1:1'b0;
assign ENABLE_NOT_G_AND_RN = (!G&RN) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_RN_AND_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_RN_AND_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_RN_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge RN, negedge G &&& (ENABLE_D_AND_SN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge RN &&& (ENABLE_NOT_G_AND_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, negedge G &&& (ENABLE_NOT_D_AND_RN == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$setuphold(posedge RN &&& (ENABLE_NOT_G == 1'b1), posedge SN, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_G_AND_RN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (Q +: 1'b0))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1)
(RN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b1)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b1 && RN==1'b0)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b0)
(negedge RN *> (QN -: 1'b0))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b1 && G==1'b1)
(RN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1 && RN==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0 && RN==1'b1)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b1 && RN==1'b0)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATSRXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATSX1 (Q, QN, D, G, SN);
output  Q, QN;
input  D, G, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_G ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_G = (!G) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, negedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_G == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && G==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATSX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATSX2 (Q, QN, D, G, SN);
output  Q, QN;
input  D, G, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_G ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_G = (!G) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, negedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_G == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && G==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATSX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATSX4 (Q, QN, D, G, SN);
output  Q, QN;
input  D, G, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_G ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_G = (!G) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, negedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_G == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && G==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATSX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATSXL (Q, QN, D, G, SN);
output  Q, QN;
input  D, G, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,G);

wire ENABLE_SN ;
wire ENABLE_NOT_D ;
wire ENABLE_NOT_G ;
assign ENABLE_SN = (SN) ? 1'b1:1'b0;
assign ENABLE_NOT_D = (!D) ? 1'b1:1'b0;
assign ENABLE_NOT_G = (!G) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_SN == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_SN == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$recrem(posedge SN, negedge G &&& (ENABLE_NOT_D == 1'b1), `ARM_RECOVERY_TIME, `ARM_REMOVAL_TIME, NOTIFIER);
$width(negedge SN &&& (ENABLE_NOT_G == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
if (D==1'b0 && G==1'b1)
(SN => Q) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge SN *> (Q +: 1'b1))=(`ARM_PROP_DELAY, `ARM_INVALID_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);
if (D==1'b0 && G==1'b1)
(SN => QN) = (`ARM_PROP_DELAY, `ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
(negedge SN *> (QN -: 1'b1))=(`ARM_INVALID_DELAY, `ARM_PROP_DELAY);

endspecify
endmodule // TLATSXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATTSCOX1 (ECKN, CKN, E, SE);
output ECKN;
input  E, SE, CKN;
reg NOTIFIER;

supply1 R, S;

  not      I0 (nclk,CKN);
  or       I1 (n1, SE, E);
  udp_tlat_PWR I2 (n0, n1, nclk, R, S, 1'b1, 1'b0, NOTIFIER);
  not      I3 (nn0,n0);
  or       I4 (ECKN, nn0, CKN);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CKN => ECKN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CKN => ECKN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CKN => ECKN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(posedge CKN => (ECKN:1'bx)) = (`ARM_PROP_DELAY,`ARM_INVALID_DELAY);
$width(posedge CKN &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(posedge CKN &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATTSCOX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATTSCOX2 (ECKN, CKN, E, SE);
output ECKN;
input  E, SE, CKN;
reg NOTIFIER;

supply1 R, S;

  not      I0 (nclk,CKN);
  or       I1 (n1, SE, E);
  udp_tlat_PWR I2 (n0, n1, nclk, R, S, 1'b1, 1'b0, NOTIFIER);
  not      I3 (nn0,n0);
  or       I4 (ECKN, nn0, CKN);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CKN => ECKN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CKN => ECKN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CKN => ECKN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(posedge CKN => (ECKN:1'bx)) = (`ARM_PROP_DELAY,`ARM_INVALID_DELAY);
$width(posedge CKN &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(posedge CKN &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATTSCOX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATTSCOX3 (ECKN, CKN, E, SE);
output ECKN;
input  E, SE, CKN;
reg NOTIFIER;

supply1 R, S;

  not      I0 (nclk,CKN);
  or       I1 (n1, SE, E);
  udp_tlat_PWR I2 (n0, n1, nclk, R, S, 1'b1, 1'b0, NOTIFIER);
  not      I3 (nn0,n0);
  or       I4 (ECKN, nn0, CKN);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CKN => ECKN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CKN => ECKN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CKN => ECKN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(posedge CKN => (ECKN:1'bx)) = (`ARM_PROP_DELAY,`ARM_INVALID_DELAY);
$width(posedge CKN &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(posedge CKN &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATTSCOX3
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATTSCOX4 (ECKN, CKN, E, SE);
output ECKN;
input  E, SE, CKN;
reg NOTIFIER;

supply1 R, S;

  not      I0 (nclk,CKN);
  or       I1 (n1, SE, E);
  udp_tlat_PWR I2 (n0, n1, nclk, R, S, 1'b1, 1'b0, NOTIFIER);
  not      I3 (nn0,n0);
  or       I4 (ECKN, nn0, CKN);


wire ENABLE_NOT_E_AND_NOT_SE ;
wire ENABLE_E_OR_SE ;
wire ENABLE_NOT_SE ;
wire ENABLE_NOT_E ;
assign ENABLE_NOT_E_AND_NOT_SE = (!E&!SE) ? 1'b1:1'b0;
assign ENABLE_E_OR_SE = (E | SE) ? 1'b1:1'b0;
assign ENABLE_NOT_SE = (!SE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;

specify
if (E==1'b0 && SE==1'b1)
(CKN => ECKN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b0)
(CKN => ECKN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b1 && SE==1'b1)
(CKN => ECKN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (E==1'b0 && SE==1'b0)
(posedge CKN => (ECKN:1'bx)) = (`ARM_PROP_DELAY,`ARM_INVALID_DELAY);
$width(posedge CKN &&& (ENABLE_NOT_E_AND_NOT_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$width(posedge CKN &&& (ENABLE_E_OR_SE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), posedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_SE == 1'b1), negedge E, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_E == 1'b1), posedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge CKN &&& (ENABLE_NOT_E == 1'b1), negedge SE, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);

endspecify
endmodule // TLATTSCOX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATX1 (Q, QN, D, G);
output  Q, QN;
input  D, G;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,G);


specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TLATX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATX2 (Q, QN, D, G);
output  Q, QN;
input  D, G;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,G);


specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TLATX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATX4 (Q, QN, D, G);
output  Q, QN;
input  D, G;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,G);


specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TLATX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TLATXL (Q, QN, D, G);
output  Q, QN;
input  D, G;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
buf      I1 (Q, n0);
not      I2 (QN, n0);
not  I3(clk,G);


specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(D => QN) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G, posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G, negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G,`ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge G => (QN:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TLATXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TTLATX1 (Q, D, G, OE);
output Q;
input  D, G, OE;
reg NOTIFIER;
supply1 RN, SN;
supply1 xRN, xSN;
supply1 dRN, dSN;

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
bufif1   I1 (Q, n0, OE);
not  I3(clk,G);

wire ENABLE_OE ;
assign ENABLE_OE = (OE) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
( OE => Q ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
( OE => Q ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (G==1'b1)
( OE => Q ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_OE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_OE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_OE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TTLATX1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TTLATX2 (Q, D, G, OE);
output Q;
input  D, G, OE;
reg NOTIFIER;
supply1 RN, SN;
supply1 xRN, xSN;
supply1 dRN, dSN;

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
bufif1   I1 (Q, n0, OE);
not  I3(clk,G);

wire ENABLE_OE ;
assign ENABLE_OE = (OE) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
( OE => Q ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
( OE => Q ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (G==1'b1)
( OE => Q ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_OE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_OE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_OE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TTLATX2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TTLATX4 (Q, D, G, OE);
output Q;
input  D, G, OE;
reg NOTIFIER;
supply1 RN, SN;
supply1 xRN, xSN;
supply1 dRN, dSN;

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
bufif1   I1 (Q, n0, OE);
not  I3(clk,G);

wire ENABLE_OE ;
assign ENABLE_OE = (OE) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
( OE => Q ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
( OE => Q ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (G==1'b1)
( OE => Q ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_OE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_OE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_OE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TTLATX4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module TTLATXL (Q, D, G, OE);
output Q;
input  D, G, OE;
reg NOTIFIER;
supply1 RN, SN;
supply1 xRN, xSN;
supply1 dRN, dSN;

udp_tlat_PWR I0 (n0, D, clk, xRN, xSN, 1'b1, 1'b0, NOTIFIER);
bufif1   I1 (Q, n0, OE);
not  I3(clk,G);

wire ENABLE_OE ;
assign ENABLE_OE = (OE) ? 1'b1:1'b0;

specify
(D => Q) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b0 && G==1'b0)
( OE => Q ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (D==1'b1 && G==1'b0)
( OE => Q ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (G==1'b1)
( OE => Q ) = (`ARM_INVALID_DELAY, `ARM_INVALID_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY,`ARM_PROP_DELAY);
$setuphold(negedge G &&& (ENABLE_OE == 1'b1), posedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$setuphold(negedge G &&& (ENABLE_OE == 1'b1), negedge D, `ARM_SETUP_TIME, `ARM_HOLD_TIME, NOTIFIER);
$width(posedge G &&& (ENABLE_OE == 1'b1), `ARM_WIDTH,`ARM_WIDTH_THD,NOTIFIER);
(posedge G => (Q:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // TTLATXL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2X1 (Y, A, B);
output Y;
input A, B;

  xnor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR2X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2X2 (Y, A, B);
output Y;
input A, B;

  xnor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR2X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2X4 (Y, A, B);
output Y;
input A, B;

  xnor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR2X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR2XL (Y, A, B);
output Y;
input A, B;

  xnor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR2XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3X2 (Y, A, B, C);
output Y;
input A, B, C;

  xnor I0(Y, A, B, C);



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR3X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XNOR3X4 (Y, A, B, C);
output Y;
input A, B, C;

  xnor I0(Y, A, B, C);



specify
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XNOR3X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2X1 (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR2X1
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2X2 (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR2X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2X4 (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR2X4
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR2XL (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);



specify
(posedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge A => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(posedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
(negedge B => (Y:1'bx)) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR2XL
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3X2 (Y, A, B, C);
output Y;
input A, B, C;

  xor I0(Y, A, B, C);



specify
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR3X2
`endcelldefine
`timescale 1ns/1ps
`celldefine
module XOR3X4 (Y, A, B, C);
output Y;
input A, B, C;

  xor I0(Y, A, B, C);



specify
if (B==1'b0 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b0 && C==1'b0)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (B==1'b1 && C==1'b1)
(A => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && C==1'b0)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && C==1'b1)
(B => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b0 && B==1'b0)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);
if (A==1'b1 && B==1'b1)
(C => Y) = (`ARM_PROP_DELAY,`ARM_PROP_DELAY);

endspecify
endmodule // XOR3X4
`endcelldefine
`endif
`endif
