////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
/// TSMC Library/IP Product
/// Filename: tcb013bcd.v
/// Technology: CM013ML,CM013MP,CV013NH,CV013NI
/// Product Type: Standard Cell
/// Product Name: tcb013bcd
/// Version: 110a
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////
///  STATEMENT OF USE
///
///  This information contains confidential and proprietary information of TSMC.
///  No part of this information may be reproduced, transmitted, transcribed,
///  stored in a retrieval system, or translated into any human or computer
///  language, in any form or by any means, electronic, mechanical, magnetic,
///  optical, chemical, manual, or otherwise, without the prior written permission
///  of TSMC.  This information was prepared for informational purpose and is for
///  use by TSMC's customers only.  TSMC reserves the right to make changes in the
///  information at any time and without notice.
///
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
`timescale 1ns/10ps

`celldefine
module AN2D0 (A1, A2, Z);
    input A1, A2;
    output Z;
    and (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN2D1 (A1, A2, Z);
    input A1, A2;
    output Z;
    and (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN2D2 (A1, A2, Z);
    input A1, A2;
    output Z;
    and (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN2D4 (A1, A2, Z);
    input A1, A2;
    output Z;
    and (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN2D8 (A1, A2, Z);
    input A1, A2;
    output Z;
    and (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN2XD1 (A1, A2, Z);
    input A1, A2;
    output Z;
    and (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN3D0 (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    and (Z, A1, A2, A3);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN3D1 (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    and (Z, A1, A2, A3);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN3D2 (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    and (Z, A1, A2, A3);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN3D4 (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    and (Z, A1, A2, A3);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN3D8 (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    and (Z, A1, A2, A3);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN3XD1 (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    and (Z, A1, A2, A3);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN4D0 (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    and (Z, A1, A2, A3, A4);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN4D1 (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    and (Z, A1, A2, A3, A4);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN4D2 (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    and (Z, A1, A2, A3, A4);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN4D4 (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    and (Z, A1, A2, A3, A4);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN4D8 (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    and (Z, A1, A2, A3, A4);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN4XD1 (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    and (Z, A1, A2, A3, A4);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ANTENNA (I);
    input I;
    buf (I_buf, I);

endmodule
`endcelldefine

`celldefine
module AO211D0 (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
    and (I0_out, A1, A2);
    or (Z, I0_out, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO211D1 (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
    and (I0_out, A1, A2);
    or (Z, I0_out, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO211D2 (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
    and (I0_out, A1, A2);
    or (Z, I0_out, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO211D4 (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
    and (I0_out, A1, A2);
    or (Z, I0_out, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO21D0 (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
    and (I0_out, A1, A2);
    or (Z, I0_out, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO21D1 (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
    and (I0_out, A1, A2);
    or (Z, I0_out, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO21D2 (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
    and (I0_out, A1, A2);
    or (Z, I0_out, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO21D4 (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
    and (I0_out, A1, A2);
    or (Z, I0_out, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO221D0 (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (Z, I0_out, I1_out, C);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO221D1 (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (Z, I0_out, I1_out, C);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO221D2 (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (Z, I0_out, I1_out, C);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO221D4 (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (Z, I0_out, I1_out, C);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO222D0 (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    and (I2_out, C1, C2);
    or (Z, I0_out, I1_out, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO222D1 (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    and (I2_out, C1, C2);
    or (Z, I0_out, I1_out, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO222D2 (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    and (I2_out, C1, C2);
    or (Z, I0_out, I1_out, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO222D4 (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    and (I2_out, C1, C2);
    or (Z, I0_out, I1_out, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO22D0 (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO22D1 (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO22D2 (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO22D4 (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO31D0 (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
    and (I0_out, A1, A2, A3);
    or (Z, I0_out, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO31D1 (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
    and (I0_out, A1, A2, A3);
    or (Z, I0_out, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO31D2 (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
    and (I0_out, A1, A2, A3);
    or (Z, I0_out, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO31D4 (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
    and (I0_out, A1, A2, A3);
    or (Z, I0_out, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO32D0 (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
    and (I0_out, A1, A2, A3);
    and (I1_out, B1, B2);
    or (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO32D1 (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
    and (I0_out, A1, A2, A3);
    and (I1_out, B1, B2);
    or (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO32D2 (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
    and (I0_out, A1, A2, A3);
    and (I1_out, B1, B2);
    or (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO32D4 (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
    and (I0_out, A1, A2, A3);
    and (I1_out, B1, B2);
    or (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO33D0 (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
    and (I0_out, A1, A2, A3);
    and (I1_out, B1, B2, B3);
    or (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO33D1 (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
    and (I0_out, A1, A2, A3);
    and (I1_out, B1, B2, B3);
    or (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO33D2 (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
    and (I0_out, A1, A2, A3);
    and (I1_out, B1, B2, B3);
    or (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO33D4 (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
    and (I0_out, A1, A2, A3);
    and (I1_out, B1, B2, B3);
    or (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI211D0 (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    and (I0_out, A1, A2);
    or (I2_out, I0_out, B, C);
    not (ZN, I2_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI211D1 (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    and (I0_out, A1, A2);
    or (I2_out, I0_out, B, C);
    not (ZN, I2_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI211D2 (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    and (I0_out, A1, A2);
    or (I2_out, I0_out, B, C);
    not (ZN, I2_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI211D4 (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    and (I0_out, A1, A2);
    or (I2_out, I0_out, B, C);
    not (ZN, I2_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI211XD0 (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    and (I0_out, A1, A2);
    or (I2_out, I0_out, B, C);
    not (ZN, I2_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI211XD1 (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    and (I0_out, A1, A2);
    or (I2_out, I0_out, B, C);
    not (ZN, I2_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI211XD2 (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    and (I0_out, A1, A2);
    or (I2_out, I0_out, B, C);
    not (ZN, I2_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI211XD4 (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    and (I0_out, A1, A2);
    or (I2_out, I0_out, B, C);
    not (ZN, I2_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI21D0 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    and (I0_out, A1, A2);
    or (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI21D1 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    and (I0_out, A1, A2);
    or (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI21D2 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    and (I0_out, A1, A2);
    or (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI21D4 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    and (I0_out, A1, A2);
    or (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI221D0 (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (I2_out, I0_out, I1_out, C);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI221D1 (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (I2_out, I0_out, I1_out, C);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI221D2 (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (I2_out, I0_out, I1_out, C);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI221D4 (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (I2_out, I0_out, I1_out, C);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI221XD4 (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (I2_out, I0_out, I1_out, C);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI222D0 (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
    and (I0_out, A1, A2);
    and (I1_out, C1, C2);
    and (I2_out, B1, B2);
    or (I3_out, I0_out, I1_out, I2_out);
    not (ZN, I3_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI222D1 (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
    and (I0_out, A1, A2);
    and (I1_out, C1, C2);
    and (I2_out, B1, B2);
    or (I3_out, I0_out, I1_out, I2_out);
    not (ZN, I3_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI222D2 (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
    and (I0_out, A1, A2);
    and (I1_out, C1, C2);
    and (I2_out, B1, B2);
    or (I3_out, I0_out, I1_out, I2_out);
    not (ZN, I3_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI222D4 (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
    and (I0_out, A1, A2);
    and (I1_out, C1, C2);
    and (I2_out, B1, B2);
    or (I3_out, I0_out, I1_out, I2_out);
    not (ZN, I3_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI222XD4 (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
    and (I0_out, A1, A2);
    and (I1_out, C1, C2);
    and (I2_out, B1, B2);
    or (I3_out, I0_out, I1_out, I2_out);
    not (ZN, I3_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI22D0 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI22D1 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI22D2 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI22D4 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI31D0 (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
    and (I0_out, A1, A2, A3);
    or (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI31D1 (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
    and (I0_out, A1, A2, A3);
    or (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI31D2 (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
    and (I0_out, A1, A2, A3);
    or (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI31D4 (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
    and (I0_out, A1, A2, A3);
    or (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI32D0 (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
    and (I0_out, B1, B2);
    and (I1_out, A1, A2, A3);
    or (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI32D1 (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
    and (I0_out, B1, B2);
    and (I1_out, A1, A2, A3);
    or (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI32D2 (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
    and (I0_out, B1, B2);
    and (I1_out, A1, A2, A3);
    or (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI32D4 (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
    and (I0_out, B1, B2);
    and (I1_out, A1, A2, A3);
    or (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI32XD4 (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
    and (I0_out, B1, B2);
    and (I1_out, A1, A2, A3);
    or (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI33D0 (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
    and (I0_out, B1, B2, B3);
    and (I1_out, A1, A2, A3);
    or (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI33D1 (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
    and (I0_out, B1, B2, B3);
    and (I1_out, A1, A2, A3);
    or (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI33D2 (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
    and (I0_out, B1, B2, B3);
    and (I1_out, A1, A2, A3);
    or (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI33D4 (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
    and (I0_out, B1, B2, B3);
    and (I1_out, A1, A2, A3);
    or (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI33XD4 (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
    and (I0_out, B1, B2, B3);
    and (I1_out, A1, A2, A3);
    or (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BENCD1 (M0, M1, M2, X2, A, S);
    input M0, M1, M2;
    output X2, A, S;
    xor (I0_out, M0, M1);
    not (X2, I0_out);
    or (I1_out, M0, M1);
    not (I2_out, I1_out);
    or (A, I2_out, M2);
    and (I3_out, M0, M1);
    not (I4_out, I3_out);
    and (I5_out, I4_out, M2);
    not (S, I5_out);

  specify
    (M0 => A) = (0, 0);
    (M1 => A) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b1)
    (M2 => A) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b0)
    (M2 => A) = (0, 0);
    if (M0 == 1'b0 && M1 == 1'b1)
    (M2 => A) = (0, 0);
    (M0 => S) = (0, 0);
    (M1 => S) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b0)
    (M2 => S) = (0, 0);
    if (M0 == 1'b0 && M1 == 1'b1)
    (M2 => S) = (0, 0);
    if (M0 == 1'b0 && M1 == 1'b0)
    (M2 => S) = (0, 0);
    if (M1 == 1'b1 && M2 == 1'b1)
    (M0 => X2) = (0, 0);
    if (M1 == 1'b1 && M2 == 1'b0)
    (M0 => X2) = (0, 0);
    if (M1 == 1'b0 && M2 == 1'b1)
    (M0 => X2) = (0, 0);
    if (M1 == 1'b0 && M2 == 1'b0)
    (M0 => X2) = (0, 0);
    if (M0 == 1'b1 && M2 == 1'b1)
    (M1 => X2) = (0, 0);
    if (M0 == 1'b1 && M2 == 1'b0)
    (M1 => X2) = (0, 0);
    if (M0 == 1'b0 && M2 == 1'b1)
    (M1 => X2) = (0, 0);
    if (M0 == 1'b0 && M2 == 1'b0)
    (M1 => X2) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BENCD2 (M0, M1, M2, X2, A, S);
    input M0, M1, M2;
    output X2, A, S;
    xor (I0_out, M0, M1);
    not (X2, I0_out);
    or (I1_out, M0, M1);
    not (I2_out, I1_out);
    or (A, I2_out, M2);
    and (I3_out, M0, M1);
    not (I4_out, I3_out);
    and (I5_out, I4_out, M2);
    not (S, I5_out);

  specify
    (M0 => A) = (0, 0);
    (M1 => A) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b1)
    (M2 => A) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b0)
    (M2 => A) = (0, 0);
    if (M0 == 1'b0 && M1 == 1'b1)
    (M2 => A) = (0, 0);
    (M0 => S) = (0, 0);
    (M1 => S) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b0)
    (M2 => S) = (0, 0);
    if (M0 == 1'b0 && M1 == 1'b1)
    (M2 => S) = (0, 0);
    if (M0 == 1'b0 && M1 == 1'b0)
    (M2 => S) = (0, 0);
    if (M1 == 1'b1 && M2 == 1'b1)
    (M0 => X2) = (0, 0);
    if (M1 == 1'b1 && M2 == 1'b0)
    (M0 => X2) = (0, 0);
    if (M1 == 1'b0 && M2 == 1'b1)
    (M0 => X2) = (0, 0);
    if (M1 == 1'b0 && M2 == 1'b0)
    (M0 => X2) = (0, 0);
    if (M0 == 1'b1 && M2 == 1'b1)
    (M1 => X2) = (0, 0);
    if (M0 == 1'b1 && M2 == 1'b0)
    (M1 => X2) = (0, 0);
    if (M0 == 1'b0 && M2 == 1'b1)
    (M1 => X2) = (0, 0);
    if (M0 == 1'b0 && M2 == 1'b0)
    (M1 => X2) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BENCD4 (M0, M1, M2, X2, A, S);
    input M0, M1, M2;
    output X2, A, S;
    xor (I0_out, M0, M1);
    not (X2, I0_out);
    or (I1_out, M0, M1);
    not (I2_out, I1_out);
    or (A, I2_out, M2);
    and (I3_out, M0, M1);
    not (I4_out, I3_out);
    and (I5_out, I4_out, M2);
    not (S, I5_out);

  specify
    (M0 => A) = (0, 0);
    (M1 => A) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b1)
    (M2 => A) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b0)
    (M2 => A) = (0, 0);
    if (M0 == 1'b0 && M1 == 1'b1)
    (M2 => A) = (0, 0);
    (M0 => S) = (0, 0);
    (M1 => S) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b0)
    (M2 => S) = (0, 0);
    if (M0 == 1'b0 && M1 == 1'b1)
    (M2 => S) = (0, 0);
    if (M0 == 1'b0 && M1 == 1'b0)
    (M2 => S) = (0, 0);
    if (M1 == 1'b1 && M2 == 1'b1)
    (M0 => X2) = (0, 0);
    if (M1 == 1'b1 && M2 == 1'b0)
    (M0 => X2) = (0, 0);
    if (M1 == 1'b0 && M2 == 1'b1)
    (M0 => X2) = (0, 0);
    if (M1 == 1'b0 && M2 == 1'b0)
    (M0 => X2) = (0, 0);
    if (M0 == 1'b1 && M2 == 1'b1)
    (M1 => X2) = (0, 0);
    if (M0 == 1'b1 && M2 == 1'b0)
    (M1 => X2) = (0, 0);
    if (M0 == 1'b0 && M2 == 1'b1)
    (M1 => X2) = (0, 0);
    if (M0 == 1'b0 && M2 == 1'b0)
    (M1 => X2) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BHD (Z);
    inout Z;
    not (weak0, weak1) (Z, Z_buf);
    not                (Z_buf, Z);

endmodule
`endcelldefine

`celldefine
module BMLD1 (X2, A, S, M0, M1, PP);
    input X2, A, S, M0, M1;
    output PP;
    tsmc_mux (I0_out, S, A, M0);
    tsmc_mux (I1_out, S, A, M1);
    tsmc_mux (I2_out, I1_out, I0_out, X2);
    not (PP, I2_out);

  specify
    if (M0 == 1'b1 && M1 == 1'b1 && S == 1'b1 && X2 == 1'b1)
    (A => PP) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b1 && S == 1'b0 && X2 == 1'b1)
    (A => PP) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b1 && S == 1'b1 && X2 == 1'b0)
    (A => PP) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b1 && S == 1'b0 && X2 == 1'b0)
    (A => PP) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b0 && S == 1'b1 && X2 == 1'b1)
    (A => PP) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b0 && S == 1'b0 && X2 == 1'b1)
    (A => PP) = (0, 0);
    if (M0 == 1'b0 && M1 == 1'b1 && S == 1'b1 && X2 == 1'b0)
    (A => PP) = (0, 0);
    if (M0 == 1'b0 && M1 == 1'b1 && S == 1'b0 && X2 == 1'b0)
    (A => PP) = (0, 0);
    if (A == 1'b0 && M1 == 1'b1 && S == 1'b1 && X2 == 1'b1)
    (M0 => PP) = (0, 0);
    if (A == 1'b0 && M1 == 1'b0 && S == 1'b1 && X2 == 1'b1)
    (M0 => PP) = (0, 0);
    if (A == 1'b1 && M1 == 1'b1 && S == 1'b0 && X2 == 1'b1)
    (M0 => PP) = (0, 0);
    if (A == 1'b1 && M1 == 1'b0 && S == 1'b0 && X2 == 1'b1)
    (M0 => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b1 && S == 1'b1 && X2 == 1'b0)
    (M1 => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b0 && S == 1'b1 && X2 == 1'b0)
    (M1 => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b1 && S == 1'b0 && X2 == 1'b0)
    (M1 => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b0 && S == 1'b0 && X2 == 1'b0)
    (M1 => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b1 && M1 == 1'b0 && X2 == 1'b0)
    (S => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b1 && M1 == 1'b0 && X2 == 1'b0)
    (S => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b0 && M1 == 1'b1 && X2 == 1'b1)
    (S => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b0 && M1 == 1'b1 && X2 == 1'b1)
    (S => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b0 && M1 == 1'b0 && X2 == 1'b1)
    (S => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b0 && M1 == 1'b0 && X2 == 1'b1)
    (S => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b0 && M1 == 1'b0 && X2 == 1'b0)
    (S => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b0 && M1 == 1'b0 && X2 == 1'b0)
    (S => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b0 && M1 == 1'b1 && S == 1'b0)
    (X2 => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b1 && M1 == 1'b0 && S == 1'b1)
    (X2 => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b1 && M1 == 1'b0 && S == 1'b0)
    (X2 => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b0 && M1 == 1'b1 && S == 1'b1)
    (X2 => PP) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BMLD2 (X2, A, S, M0, M1, PP);
    input X2, A, S, M0, M1;
    output PP;
    tsmc_mux (I0_out, S, A, M0);
    tsmc_mux (I1_out, S, A, M1);
    tsmc_mux (I2_out, I1_out, I0_out, X2);
    not (PP, I2_out);

  specify
    if (M0 == 1'b1 && M1 == 1'b1 && S == 1'b1 && X2 == 1'b1)
    (A => PP) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b1 && S == 1'b0 && X2 == 1'b1)
    (A => PP) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b1 && S == 1'b1 && X2 == 1'b0)
    (A => PP) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b1 && S == 1'b0 && X2 == 1'b0)
    (A => PP) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b0 && S == 1'b1 && X2 == 1'b1)
    (A => PP) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b0 && S == 1'b0 && X2 == 1'b1)
    (A => PP) = (0, 0);
    if (M0 == 1'b0 && M1 == 1'b1 && S == 1'b1 && X2 == 1'b0)
    (A => PP) = (0, 0);
    if (M0 == 1'b0 && M1 == 1'b1 && S == 1'b0 && X2 == 1'b0)
    (A => PP) = (0, 0);
    if (A == 1'b0 && M1 == 1'b1 && S == 1'b1 && X2 == 1'b1)
    (M0 => PP) = (0, 0);
    if (A == 1'b0 && M1 == 1'b0 && S == 1'b1 && X2 == 1'b1)
    (M0 => PP) = (0, 0);
    if (A == 1'b1 && M1 == 1'b1 && S == 1'b0 && X2 == 1'b1)
    (M0 => PP) = (0, 0);
    if (A == 1'b1 && M1 == 1'b0 && S == 1'b0 && X2 == 1'b1)
    (M0 => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b1 && S == 1'b1 && X2 == 1'b0)
    (M1 => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b0 && S == 1'b1 && X2 == 1'b0)
    (M1 => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b1 && S == 1'b0 && X2 == 1'b0)
    (M1 => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b0 && S == 1'b0 && X2 == 1'b0)
    (M1 => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b1 && M1 == 1'b0 && X2 == 1'b0)
    (S => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b1 && M1 == 1'b0 && X2 == 1'b0)
    (S => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b0 && M1 == 1'b1 && X2 == 1'b1)
    (S => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b0 && M1 == 1'b1 && X2 == 1'b1)
    (S => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b0 && M1 == 1'b0 && X2 == 1'b1)
    (S => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b0 && M1 == 1'b0 && X2 == 1'b1)
    (S => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b0 && M1 == 1'b0 && X2 == 1'b0)
    (S => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b0 && M1 == 1'b0 && X2 == 1'b0)
    (S => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b0 && M1 == 1'b1 && S == 1'b0)
    (X2 => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b1 && M1 == 1'b0 && S == 1'b1)
    (X2 => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b1 && M1 == 1'b0 && S == 1'b0)
    (X2 => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b0 && M1 == 1'b1 && S == 1'b1)
    (X2 => PP) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BMLD4 (X2, A, S, M0, M1, PP);
    input X2, A, S, M0, M1;
    output PP;
    tsmc_mux (I0_out, S, A, M0);
    tsmc_mux (I1_out, S, A, M1);
    tsmc_mux (I2_out, I1_out, I0_out, X2);
    not (PP, I2_out);

  specify
    if (M0 == 1'b1 && M1 == 1'b1 && S == 1'b1 && X2 == 1'b1)
    (A => PP) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b1 && S == 1'b0 && X2 == 1'b1)
    (A => PP) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b1 && S == 1'b1 && X2 == 1'b0)
    (A => PP) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b1 && S == 1'b0 && X2 == 1'b0)
    (A => PP) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b0 && S == 1'b1 && X2 == 1'b1)
    (A => PP) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b0 && S == 1'b0 && X2 == 1'b1)
    (A => PP) = (0, 0);
    if (M0 == 1'b0 && M1 == 1'b1 && S == 1'b1 && X2 == 1'b0)
    (A => PP) = (0, 0);
    if (M0 == 1'b0 && M1 == 1'b1 && S == 1'b0 && X2 == 1'b0)
    (A => PP) = (0, 0);
    if (A == 1'b0 && M1 == 1'b1 && S == 1'b1 && X2 == 1'b1)
    (M0 => PP) = (0, 0);
    if (A == 1'b0 && M1 == 1'b0 && S == 1'b1 && X2 == 1'b1)
    (M0 => PP) = (0, 0);
    if (A == 1'b1 && M1 == 1'b1 && S == 1'b0 && X2 == 1'b1)
    (M0 => PP) = (0, 0);
    if (A == 1'b1 && M1 == 1'b0 && S == 1'b0 && X2 == 1'b1)
    (M0 => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b1 && S == 1'b1 && X2 == 1'b0)
    (M1 => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b0 && S == 1'b1 && X2 == 1'b0)
    (M1 => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b1 && S == 1'b0 && X2 == 1'b0)
    (M1 => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b0 && S == 1'b0 && X2 == 1'b0)
    (M1 => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b1 && M1 == 1'b0 && X2 == 1'b0)
    (S => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b1 && M1 == 1'b0 && X2 == 1'b0)
    (S => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b0 && M1 == 1'b1 && X2 == 1'b1)
    (S => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b0 && M1 == 1'b1 && X2 == 1'b1)
    (S => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b0 && M1 == 1'b0 && X2 == 1'b1)
    (S => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b0 && M1 == 1'b0 && X2 == 1'b1)
    (S => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b0 && M1 == 1'b0 && X2 == 1'b0)
    (S => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b0 && M1 == 1'b0 && X2 == 1'b0)
    (S => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b0 && M1 == 1'b1 && S == 1'b0)
    (X2 => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b1 && M1 == 1'b0 && S == 1'b1)
    (X2 => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b1 && M1 == 1'b0 && S == 1'b0)
    (X2 => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b0 && M1 == 1'b1 && S == 1'b1)
    (X2 => PP) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFFD0 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFFD1 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFFD12 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFFD16 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFFD2 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFFD20 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFFD24 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFFD3 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFFD4 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFFD6 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFFD8 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFTD0 (I, OE, Z);
    input I, OE;
    output Z;
    bufif1 (Z, I, OE);

  specify
    (I => Z) = (0, 0);
    (OE => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFTD1 (I, OE, Z);
    input I, OE;
    output Z;
    bufif1 (Z, I, OE);

  specify
    (I => Z) = (0, 0);
    (OE => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFTD12 (I, OE, Z);
    input I, OE;
    output Z;
    bufif1 (Z, I, OE);

  specify
    (I => Z) = (0, 0);
    (OE => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFTD16 (I, OE, Z);
    input I, OE;
    output Z;
    bufif1 (Z, I, OE);

  specify
    (I => Z) = (0, 0);
    (OE => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFTD2 (I, OE, Z);
    input I, OE;
    output Z;
    bufif1 (Z, I, OE);

  specify
    (I => Z) = (0, 0);
    (OE => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFTD20 (I, OE, Z);
    input I, OE;
    output Z;
    bufif1 (Z, I, OE);

  specify
    (I => Z) = (0, 0);
    (OE => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFTD24 (I, OE, Z);
    input I, OE;
    output Z;
    bufif1 (Z, I, OE);

  specify
    (I => Z) = (0, 0);
    (OE => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFTD3 (I, OE, Z);
    input I, OE;
    output Z;
    bufif1 (Z, I, OE);

  specify
    (I => Z) = (0, 0);
    (OE => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFTD4 (I, OE, Z);
    input I, OE;
    output Z;
    bufif1 (Z, I, OE);

  specify
    (I => Z) = (0, 0);
    (OE => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFTD6 (I, OE, Z);
    input I, OE;
    output Z;
    bufif1 (Z, I, OE);

  specify
    (I => Z) = (0, 0);
    (OE => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFTD8 (I, OE, Z);
    input I, OE;
    output Z;
    bufif1 (Z, I, OE);

  specify
    (I => Z) = (0, 0);
    (OE => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKAN2D0 (A1, A2, Z);
    input A1, A2;
    output Z;
    and (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKAN2D1 (A1, A2, Z);
    input A1, A2;
    output Z;
    and (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKAN2D2 (A1, A2, Z);
    input A1, A2;
    output Z;
    and (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKAN2D4 (A1, A2, Z);
    input A1, A2;
    output Z;
    and (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKAN2D8 (A1, A2, Z);
    input A1, A2;
    output Z;
    and (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBD0 (CLK, C);
    input CLK;
    output C;
    buf (C, CLK);

  specify
    (CLK => C) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBD1 (CLK, C);
    input CLK;
    output C;
    buf (C, CLK);

  specify
    (CLK => C) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBD12 (CLK, C);
    input CLK;
    output C;
    buf (C, CLK);

  specify
    (CLK => C) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBD16 (CLK, C);
    input CLK;
    output C;
    buf (C, CLK);

  specify
    (CLK => C) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBD2 (CLK, C);
    input CLK;
    output C;
    buf (C, CLK);

  specify
    (CLK => C) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBD20 (CLK, C);
    input CLK;
    output C;
    buf (C, CLK);

  specify
    (CLK => C) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBD24 (CLK, C);
    input CLK;
    output C;
    buf (C, CLK);

  specify
    (CLK => C) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBD3 (CLK, C);
    input CLK;
    output C;
    buf (C, CLK);

  specify
    (CLK => C) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBD4 (CLK, C);
    input CLK;
    output C;
    buf (C, CLK);

  specify
    (CLK => C) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBD6 (CLK, C);
    input CLK;
    output C;
    buf (C, CLK);

  specify
    (CLK => C) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBD8 (CLK, C);
    input CLK;
    output C;
    buf (C, CLK);

  specify
    (CLK => C) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBXD0 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBXD1 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBXD12 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBXD16 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBXD2 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBXD20 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBXD24 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBXD3 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBXD4 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBXD6 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBXD8 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKLHQD1 ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, CPN_d, E_d;
        buf (_TE, TE_d);
        buf (_CPN, CPN_d);
        buf (_E, E_d);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `else 
        buf (_TE, TE);
        buf (_CPN, CPN);
        buf (_E, E);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
  `endif

    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (E == 1'b0 && TE == 1'b0)
    (posedge CPN => (Q+:1'b1)) = (0, 0);
    if (E == 1'b1 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CPN => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    $width (posedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CPN_d, TE_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CPN_d, TE_d);
  `else
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLHQD12 ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, CPN_d, E_d;
        buf (_TE, TE_d);
        buf (_CPN, CPN_d);
        buf (_E, E_d);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `else 
        buf (_TE, TE);
        buf (_CPN, CPN);
        buf (_E, E);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
  `endif

    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (E == 1'b0 && TE == 1'b0)
    (posedge CPN => (Q+:1'b1)) = (0, 0);
    if (E == 1'b1 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CPN => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    $width (posedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CPN_d, TE_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CPN_d, TE_d);
  `else
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLHQD16 ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, CPN_d, E_d;
        buf (_TE, TE_d);
        buf (_CPN, CPN_d);
        buf (_E, E_d);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `else 
        buf (_TE, TE);
        buf (_CPN, CPN);
        buf (_E, E);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
  `endif

    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (E == 1'b0 && TE == 1'b0)
    (posedge CPN => (Q+:1'b1)) = (0, 0);
    if (E == 1'b1 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CPN => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    $width (posedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CPN_d, TE_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CPN_d, TE_d);
  `else
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLHQD2 ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, CPN_d, E_d;
        buf (_TE, TE_d);
        buf (_CPN, CPN_d);
        buf (_E, E_d);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `else 
        buf (_TE, TE);
        buf (_CPN, CPN);
        buf (_E, E);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
  `endif

    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (E == 1'b0 && TE == 1'b0)
    (posedge CPN => (Q+:1'b1)) = (0, 0);
    if (E == 1'b1 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CPN => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    $width (posedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CPN_d, TE_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CPN_d, TE_d);
  `else
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLHQD20 ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, CPN_d, E_d;
        buf (_TE, TE_d);
        buf (_CPN, CPN_d);
        buf (_E, E_d);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `else 
        buf (_TE, TE);
        buf (_CPN, CPN);
        buf (_E, E);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
  `endif

    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (E == 1'b0 && TE == 1'b0)
    (posedge CPN => (Q+:1'b1)) = (0, 0);
    if (E == 1'b1 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CPN => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    $width (posedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CPN_d, TE_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CPN_d, TE_d);
  `else
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLHQD24 ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, CPN_d, E_d;
        buf (_TE, TE_d);
        buf (_CPN, CPN_d);
        buf (_E, E_d);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `else 
        buf (_TE, TE);
        buf (_CPN, CPN);
        buf (_E, E);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
  `endif

    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (E == 1'b0 && TE == 1'b0)
    (posedge CPN => (Q+:1'b1)) = (0, 0);
    if (E == 1'b1 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CPN => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    $width (posedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CPN_d, TE_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CPN_d, TE_d);
  `else
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLHQD3 ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, CPN_d, E_d;
        buf (_TE, TE_d);
        buf (_CPN, CPN_d);
        buf (_E, E_d);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `else 
        buf (_TE, TE);
        buf (_CPN, CPN);
        buf (_E, E);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
  `endif

    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (E == 1'b0 && TE == 1'b0)
    (posedge CPN => (Q+:1'b1)) = (0, 0);
    if (E == 1'b1 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CPN => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    $width (posedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CPN_d, TE_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CPN_d, TE_d);
  `else
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLHQD4 ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, CPN_d, E_d;
        buf (_TE, TE_d);
        buf (_CPN, CPN_d);
        buf (_E, E_d);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `else 
        buf (_TE, TE);
        buf (_CPN, CPN);
        buf (_E, E);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
  `endif

    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (E == 1'b0 && TE == 1'b0)
    (posedge CPN => (Q+:1'b1)) = (0, 0);
    if (E == 1'b1 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CPN => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    $width (posedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CPN_d, TE_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CPN_d, TE_d);
  `else
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLHQD6 ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, CPN_d, E_d;
        buf (_TE, TE_d);
        buf (_CPN, CPN_d);
        buf (_E, E_d);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `else 
        buf (_TE, TE);
        buf (_CPN, CPN);
        buf (_E, E);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
  `endif

    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (E == 1'b0 && TE == 1'b0)
    (posedge CPN => (Q+:1'b1)) = (0, 0);
    if (E == 1'b1 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CPN => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    $width (posedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CPN_d, TE_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CPN_d, TE_d);
  `else
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLHQD8 ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, CPN_d, E_d;
        buf (_TE, TE_d);
        buf (_CPN, CPN_d);
        buf (_E, E_d);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `else 
        buf (_TE, TE);
        buf (_CPN, CPN);
        buf (_E, E);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
  `endif

    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (E == 1'b0 && TE == 1'b0)
    (posedge CPN => (Q+:1'b1)) = (0, 0);
    if (E == 1'b1 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CPN => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    $width (posedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CPN_d, TE_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CPN_d, TE_d);
  `else
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLNQD1 (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, E_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        or (D_i, E_d, TE_d);
        not (CPB, CP_d);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP_d);
    `else 
        pullup (CDN);
        pullup (SDN);
        or (D_i, E, TE);
        not (CPB, CP);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
  `endif

    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (E == 1'b1 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b0)
    (negedge CP => (Q+:1'b0)) = (0, 0);
    $width (posedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CP_d, TE_d);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CP_d, TE_d);
  `else
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLNQD12 (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, E_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        or (D_i, E_d, TE_d);
        not (CPB, CP_d);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP_d);
    `else 
        pullup (CDN);
        pullup (SDN);
        or (D_i, E, TE);
        not (CPB, CP);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
  `endif

    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (E == 1'b1 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b0)
    (negedge CP => (Q+:1'b0)) = (0, 0);
    $width (posedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CP_d, TE_d);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CP_d, TE_d);
  `else
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLNQD16 (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, E_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        or (D_i, E_d, TE_d);
        not (CPB, CP_d);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP_d);
    `else 
        pullup (CDN);
        pullup (SDN);
        or (D_i, E, TE);
        not (CPB, CP);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
  `endif

    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (E == 1'b1 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b0)
    (negedge CP => (Q+:1'b0)) = (0, 0);
    $width (posedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CP_d, TE_d);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CP_d, TE_d);
  `else
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLNQD2 (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, E_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        or (D_i, E_d, TE_d);
        not (CPB, CP_d);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP_d);
    `else 
        pullup (CDN);
        pullup (SDN);
        or (D_i, E, TE);
        not (CPB, CP);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
  `endif

    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (E == 1'b1 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b0)
    (negedge CP => (Q+:1'b0)) = (0, 0);
    $width (posedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CP_d, TE_d);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CP_d, TE_d);
  `else
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLNQD20 (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, E_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        or (D_i, E_d, TE_d);
        not (CPB, CP_d);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP_d);
    `else 
        pullup (CDN);
        pullup (SDN);
        or (D_i, E, TE);
        not (CPB, CP);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
  `endif

    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (E == 1'b1 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b0)
    (negedge CP => (Q+:1'b0)) = (0, 0);
    $width (posedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CP_d, TE_d);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CP_d, TE_d);
  `else
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLNQD24 (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, E_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        or (D_i, E_d, TE_d);
        not (CPB, CP_d);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP_d);
    `else 
        pullup (CDN);
        pullup (SDN);
        or (D_i, E, TE);
        not (CPB, CP);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
  `endif

    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (E == 1'b1 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b0)
    (negedge CP => (Q+:1'b0)) = (0, 0);
    $width (posedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CP_d, TE_d);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CP_d, TE_d);
  `else
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLNQD3 (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, E_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        or (D_i, E_d, TE_d);
        not (CPB, CP_d);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP_d);
    `else 
        pullup (CDN);
        pullup (SDN);
        or (D_i, E, TE);
        not (CPB, CP);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
  `endif

    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (E == 1'b1 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b0)
    (negedge CP => (Q+:1'b0)) = (0, 0);
    $width (posedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CP_d, TE_d);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CP_d, TE_d);
  `else
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLNQD4 (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, E_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        or (D_i, E_d, TE_d);
        not (CPB, CP_d);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP_d);
    `else 
        pullup (CDN);
        pullup (SDN);
        or (D_i, E, TE);
        not (CPB, CP);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
  `endif

    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (E == 1'b1 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b0)
    (negedge CP => (Q+:1'b0)) = (0, 0);
    $width (posedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CP_d, TE_d);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CP_d, TE_d);
  `else
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLNQD6 (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, E_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        or (D_i, E_d, TE_d);
        not (CPB, CP_d);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP_d);
    `else 
        pullup (CDN);
        pullup (SDN);
        or (D_i, E, TE);
        not (CPB, CP);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
  `endif

    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (E == 1'b1 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b0)
    (negedge CP => (Q+:1'b0)) = (0, 0);
    $width (posedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CP_d, TE_d);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CP_d, TE_d);
  `else
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLNQD8 (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, E_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        or (D_i, E_d, TE_d);
        not (CPB, CP_d);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP_d);
    `else 
        pullup (CDN);
        pullup (SDN);
        or (D_i, E, TE);
        not (CPB, CP);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
  `endif

    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (E == 1'b1 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b0)
    (negedge CP => (Q+:1'b0)) = (0, 0);
    $width (posedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CP_d, TE_d);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CP_d, TE_d);
  `else
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKMUX2D0 (I0, I1, S, Z);
    input I0, I1, S;
    output Z;
    tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKMUX2D1 (I0, I1, S, Z);
    input I0, I1, S;
    output Z;
    tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKMUX2D2 (I0, I1, S, Z);
    input I0, I1, S;
    output Z;
    tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKMUX2D4 (I0, I1, S, Z);
    input I0, I1, S;
    output Z;
    tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND0 (CLK, CN);
    input CLK;
    output CN;
    not (CN, CLK);

  specify
    (CLK => CN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND1 (CLK, CN);
    input CLK;
    output CN;
    not (CN, CLK);

  specify
    (CLK => CN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND12 (CLK, CN);
    input CLK;
    output CN;
    not (CN, CLK);

  specify
    (CLK => CN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND16 (CLK, CN);
    input CLK;
    output CN;
    not (CN, CLK);

  specify
    (CLK => CN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND2 (CLK, CN);
    input CLK;
    output CN;
    not (CN, CLK);

  specify
    (CLK => CN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND20 (CLK, CN);
    input CLK;
    output CN;
    not (CN, CLK);

  specify
    (CLK => CN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND24 (CLK, CN);
    input CLK;
    output CN;
    not (CN, CLK);

  specify
    (CLK => CN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND2D0 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND2D1 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND2D2 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND2D3 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND2D4 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND2D8 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND3 (CLK, CN);
    input CLK;
    output CN;
    not (CN, CLK);

  specify
    (CLK => CN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND4 (CLK, CN);
    input CLK;
    output CN;
    not (CN, CLK);

  specify
    (CLK => CN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND6 (CLK, CN);
    input CLK;
    output CN;
    not (CN, CLK);

  specify
    (CLK => CN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND8 (CLK, CN);
    input CLK;
    output CN;
    not (CN, CLK);

  specify
    (CLK => CN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKNXD0 (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKNXD1 (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKNXD12 (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKNXD16 (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKNXD2 (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKNXD20 (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKNXD24 (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKNXD3 (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKNXD4 (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKNXD6 (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKNXD8 (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKXOR2D0 (A1, A2, Z);
    input A1, A2;
    output Z;
    xor (Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKXOR2D1 (A1, A2, Z);
    input A1, A2;
    output Z;
    xor (Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKXOR2D2 (A1, A2, Z);
    input A1, A2;
    output Z;
    xor (Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKXOR2D4 (A1, A2, Z);
    input A1, A2;
    output Z;
    xor (Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CMPE22D1 (A, B, S, CO);
input A, B;
output S, CO;
  xor (S, A, B);
  and (CO, A, B);

  specify
    (A => CO) = (0, 0);
    (B => CO) = (0, 0);
    if (B == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1)
    (B => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CMPE22D2 (A, B, S, CO);
input A, B;
output S, CO;
  xor (S, A, B);
  and (CO, A, B);

  specify
    (A => CO) = (0, 0);
    (B => CO) = (0, 0);
    if (B == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1)
    (B => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CMPE32D1 (A, B, CI, S, CO);
input A, B, CI;
output S, CO;
  xor  (I0_out, A, B);
  xor  (S, I0_out, CI);
  and  (I1_out, A, B);
  and  (I2_out, A, CI);
  and  (I3_out, B, CI);
  or   (CO, I1_out, I2_out, I3_out);

  specify
    if (B == 1'b1 && CI == 1'b0)
    (A => CO) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => CO) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => CO) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => CO) = (0, 0);
    if (B == 1'b1 && CI == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1)
    (CI => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CMPE32D2 (A, B, CI, S, CO);
input A, B, CI;
output S, CO;
  xor  (I0_out, A, B);
  xor  (S, I0_out, CI);
  and  (I1_out, A, B);
  and  (I2_out, A, CI);
  and  (I3_out, B, CI);
  or   (CO, I1_out, I2_out, I3_out);

  specify
    if (B == 1'b1 && CI == 1'b0)
    (A => CO) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => CO) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => CO) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => CO) = (0, 0);
    if (B == 1'b1 && CI == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1)
    (CI => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CMPE42D1 (A, B, C, D, CIX, S, COX, CO);
    input A, B, C, D, CIX;
    output S, COX, CO;
    xor (I0_out, A, B);
    xor (I1_out, I0_out, C);
    xor (I2_out, I1_out, CIX);
    xor (S, I2_out, D);
    xor (I3_out, A, B);
    xor (I4_out, I3_out, C);
    and (I5_out, I4_out, CIX);
    and (I6_out, CIX, D);
    xor (I7_out, A, B);
    xor (I8_out, I7_out, C);
    and (I9_out, I8_out, D);
    or (CO, I5_out, I6_out, I9_out);
    and (I10_out, A, B);
    and (I11_out, B, C);
    and (I12_out, A, C);
    or (COX, I10_out, I11_out, I12_out);

  specify
    if (B == 1'b1 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (A => CO) = (0, 0);
    if (B == 1'b1 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (A => CO) = (0, 0);
    if (B == 1'b0 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (A => CO) = (0, 0);
    if (B == 1'b0 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (A => CO) = (0, 0);
    if (B == 1'b1 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (A => CO) = (0, 0);
    if (B == 1'b1 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (A => CO) = (0, 0);
    if (B == 1'b0 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (A => CO) = (0, 0);
    if (B == 1'b0 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (A => CO) = (0, 0);
    if (A == 1'b1 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (B => CO) = (0, 0);
    if (A == 1'b1 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b0 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (B => CO) = (0, 0);
    if (A == 1'b0 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b1 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (B => CO) = (0, 0);
    if (A == 1'b1 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b0 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (B => CO) = (0, 0);
    if (A == 1'b0 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (C => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (C => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (C => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (C => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (C => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (C => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (C => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (C => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0)
    (CIX => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b0 && D == 1'b1)
    (CIX => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b1)
    (CIX => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0)
    (CIX => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b1)
    (CIX => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b0)
    (CIX => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b1 && D == 1'b0)
    (CIX => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b1)
    (CIX => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b1 && CIX == 1'b0)
    (D => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b1 && CIX == 1'b0)
    (D => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b0 && CIX == 1'b1)
    (D => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b0 && CIX == 1'b1)
    (D => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b1 && CIX == 1'b1)
    (D => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b1 && CIX == 1'b1)
    (D => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b0 && CIX == 1'b0)
    (D => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b0 && CIX == 1'b0)
    (D => CO) = (0, 0);
    if (B == 1'b1 && C == 1'b0 && CIX == 1'b1 && D == 1'b1)
    (A => COX) = (0, 0);
    if (B == 1'b1 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (A => COX) = (0, 0);
    if (B == 1'b1 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (A => COX) = (0, 0);
    if (B == 1'b1 && C == 1'b0 && CIX == 1'b0 && D == 1'b0)
    (A => COX) = (0, 0);
    if (B == 1'b0 && C == 1'b1 && CIX == 1'b1 && D == 1'b1)
    (A => COX) = (0, 0);
    if (B == 1'b0 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (A => COX) = (0, 0);
    if (B == 1'b0 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (A => COX) = (0, 0);
    if (B == 1'b0 && C == 1'b1 && CIX == 1'b0 && D == 1'b0)
    (A => COX) = (0, 0);
    if (A == 1'b1 && C == 1'b0 && CIX == 1'b1 && D == 1'b1)
    (B => COX) = (0, 0);
    if (A == 1'b1 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (B => COX) = (0, 0);
    if (A == 1'b1 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (B => COX) = (0, 0);
    if (A == 1'b1 && C == 1'b0 && CIX == 1'b0 && D == 1'b0)
    (B => COX) = (0, 0);
    if (A == 1'b0 && C == 1'b1 && CIX == 1'b1 && D == 1'b1)
    (B => COX) = (0, 0);
    if (A == 1'b0 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (B => COX) = (0, 0);
    if (A == 1'b0 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (B => COX) = (0, 0);
    if (A == 1'b0 && C == 1'b1 && CIX == 1'b0 && D == 1'b0)
    (B => COX) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIX == 1'b1 && D == 1'b1)
    (C => COX) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIX == 1'b1 && D == 1'b1)
    (C => COX) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (C => COX) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (C => COX) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (C => COX) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (C => COX) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIX == 1'b0 && D == 1'b0)
    (C => COX) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIX == 1'b0 && D == 1'b0)
    (C => COX) = (0, 0);
    if (B == 1'b1 && C == 1'b1 && CIX == 1'b1 && D == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && C == 1'b1 && CIX == 1'b0 && D == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && C == 1'b0 && CIX == 1'b1 && D == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && C == 1'b0 && CIX == 1'b0 && D == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && C == 1'b0 && CIX == 1'b1 && D == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && C == 1'b0 && CIX == 1'b0 && D == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && C == 1'b1 && CIX == 1'b1 && D == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && C == 1'b1 && CIX == 1'b0 && D == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b1 && C == 1'b1 && CIX == 1'b1 && D == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && C == 1'b1 && CIX == 1'b0 && D == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && C == 1'b0 && CIX == 1'b1 && D == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && C == 1'b0 && CIX == 1'b0 && D == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && C == 1'b0 && CIX == 1'b1 && D == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && C == 1'b0 && CIX == 1'b0 && D == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && C == 1'b1 && CIX == 1'b1 && D == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && C == 1'b1 && CIX == 1'b0 && D == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIX == 1'b1 && D == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIX == 1'b1 && D == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIX == 1'b0 && D == 1'b0)
    (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIX == 1'b0 && D == 1'b0)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIX == 1'b1 && D == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIX == 1'b1 && D == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIX == 1'b0 && D == 1'b0)
    (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIX == 1'b0 && D == 1'b0)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b1)
    (CIX => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b0 && D == 1'b0)
    (CIX => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
    (CIX => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
    (CIX => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
    (CIX => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
    (CIX => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b1 && D == 1'b1)
    (CIX => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b0)
    (CIX => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0)
    (CIX => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b0 && D == 1'b1)
    (CIX => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b1)
    (CIX => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0)
    (CIX => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b1)
    (CIX => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b0)
    (CIX => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b1 && D == 1'b0)
    (CIX => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b1)
    (CIX => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b1 && CIX == 1'b1)
    (D => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b1 && CIX == 1'b1)
    (D => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b0 && CIX == 1'b0)
    (D => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b0 && CIX == 1'b0)
    (D => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b1 && CIX == 1'b0)
    (D => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b1 && CIX == 1'b0)
    (D => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b0 && CIX == 1'b1)
    (D => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b0 && CIX == 1'b1)
    (D => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b1 && CIX == 1'b0)
    (D => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b1 && CIX == 1'b0)
    (D => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b0 && CIX == 1'b1)
    (D => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b0 && CIX == 1'b1)
    (D => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b1 && CIX == 1'b1)
    (D => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b1 && CIX == 1'b1)
    (D => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b0 && CIX == 1'b0)
    (D => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b0 && CIX == 1'b0)
    (D => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CMPE42D2 (A, B, C, D, CIX, S, COX, CO);
    input A, B, C, D, CIX;
    output S, COX, CO;
    xor (I0_out, A, B);
    xor (I1_out, I0_out, C);
    xor (I2_out, I1_out, CIX);
    xor (S, I2_out, D);
    xor (I3_out, A, B);
    xor (I4_out, I3_out, C);
    and (I5_out, I4_out, CIX);
    and (I6_out, CIX, D);
    xor (I7_out, A, B);
    xor (I8_out, I7_out, C);
    and (I9_out, I8_out, D);
    or (CO, I5_out, I6_out, I9_out);
    and (I10_out, A, B);
    and (I11_out, B, C);
    and (I12_out, A, C);
    or (COX, I10_out, I11_out, I12_out);

  specify
    if (B == 1'b1 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (A => CO) = (0, 0);
    if (B == 1'b1 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (A => CO) = (0, 0);
    if (B == 1'b0 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (A => CO) = (0, 0);
    if (B == 1'b0 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (A => CO) = (0, 0);
    if (B == 1'b1 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (A => CO) = (0, 0);
    if (B == 1'b1 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (A => CO) = (0, 0);
    if (B == 1'b0 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (A => CO) = (0, 0);
    if (B == 1'b0 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (A => CO) = (0, 0);
    if (A == 1'b1 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (B => CO) = (0, 0);
    if (A == 1'b1 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b0 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (B => CO) = (0, 0);
    if (A == 1'b0 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b1 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (B => CO) = (0, 0);
    if (A == 1'b1 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b0 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (B => CO) = (0, 0);
    if (A == 1'b0 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (C => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (C => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (C => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (C => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (C => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (C => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (C => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (C => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0)
    (CIX => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b0 && D == 1'b1)
    (CIX => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b1)
    (CIX => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0)
    (CIX => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b1)
    (CIX => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b0)
    (CIX => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b1 && D == 1'b0)
    (CIX => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b1)
    (CIX => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b1 && CIX == 1'b0)
    (D => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b1 && CIX == 1'b0)
    (D => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b0 && CIX == 1'b1)
    (D => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b0 && CIX == 1'b1)
    (D => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b1 && CIX == 1'b1)
    (D => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b1 && CIX == 1'b1)
    (D => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b0 && CIX == 1'b0)
    (D => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b0 && CIX == 1'b0)
    (D => CO) = (0, 0);
    if (B == 1'b1 && C == 1'b0 && CIX == 1'b1 && D == 1'b1)
    (A => COX) = (0, 0);
    if (B == 1'b1 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (A => COX) = (0, 0);
    if (B == 1'b1 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (A => COX) = (0, 0);
    if (B == 1'b1 && C == 1'b0 && CIX == 1'b0 && D == 1'b0)
    (A => COX) = (0, 0);
    if (B == 1'b0 && C == 1'b1 && CIX == 1'b1 && D == 1'b1)
    (A => COX) = (0, 0);
    if (B == 1'b0 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (A => COX) = (0, 0);
    if (B == 1'b0 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (A => COX) = (0, 0);
    if (B == 1'b0 && C == 1'b1 && CIX == 1'b0 && D == 1'b0)
    (A => COX) = (0, 0);
    if (A == 1'b1 && C == 1'b0 && CIX == 1'b1 && D == 1'b1)
    (B => COX) = (0, 0);
    if (A == 1'b1 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (B => COX) = (0, 0);
    if (A == 1'b1 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (B => COX) = (0, 0);
    if (A == 1'b1 && C == 1'b0 && CIX == 1'b0 && D == 1'b0)
    (B => COX) = (0, 0);
    if (A == 1'b0 && C == 1'b1 && CIX == 1'b1 && D == 1'b1)
    (B => COX) = (0, 0);
    if (A == 1'b0 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (B => COX) = (0, 0);
    if (A == 1'b0 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (B => COX) = (0, 0);
    if (A == 1'b0 && C == 1'b1 && CIX == 1'b0 && D == 1'b0)
    (B => COX) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIX == 1'b1 && D == 1'b1)
    (C => COX) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIX == 1'b1 && D == 1'b1)
    (C => COX) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (C => COX) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (C => COX) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (C => COX) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (C => COX) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIX == 1'b0 && D == 1'b0)
    (C => COX) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIX == 1'b0 && D == 1'b0)
    (C => COX) = (0, 0);
    if (B == 1'b1 && C == 1'b1 && CIX == 1'b1 && D == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && C == 1'b1 && CIX == 1'b0 && D == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && C == 1'b0 && CIX == 1'b1 && D == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && C == 1'b0 && CIX == 1'b0 && D == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && C == 1'b0 && CIX == 1'b1 && D == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && C == 1'b0 && CIX == 1'b0 && D == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && C == 1'b1 && CIX == 1'b1 && D == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && C == 1'b1 && CIX == 1'b0 && D == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b1 && C == 1'b1 && CIX == 1'b1 && D == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && C == 1'b1 && CIX == 1'b0 && D == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && C == 1'b0 && CIX == 1'b1 && D == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && C == 1'b0 && CIX == 1'b0 && D == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && C == 1'b0 && CIX == 1'b1 && D == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && C == 1'b0 && CIX == 1'b0 && D == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && C == 1'b1 && CIX == 1'b1 && D == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && C == 1'b1 && CIX == 1'b0 && D == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIX == 1'b1 && D == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIX == 1'b1 && D == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIX == 1'b0 && D == 1'b0)
    (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIX == 1'b0 && D == 1'b0)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIX == 1'b1 && D == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIX == 1'b1 && D == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIX == 1'b0 && D == 1'b0)
    (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIX == 1'b0 && D == 1'b0)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b1)
    (CIX => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b0 && D == 1'b0)
    (CIX => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b0)
    (CIX => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b1)
    (CIX => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b0)
    (CIX => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b1)
    (CIX => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b1 && D == 1'b1)
    (CIX => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b0)
    (CIX => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0)
    (CIX => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b0 && D == 1'b1)
    (CIX => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b1)
    (CIX => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0)
    (CIX => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b1)
    (CIX => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b0)
    (CIX => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b1 && D == 1'b0)
    (CIX => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b1)
    (CIX => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b1 && CIX == 1'b1)
    (D => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b1 && CIX == 1'b1)
    (D => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b0 && CIX == 1'b0)
    (D => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b0 && CIX == 1'b0)
    (D => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b1 && CIX == 1'b0)
    (D => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b1 && CIX == 1'b0)
    (D => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b0 && CIX == 1'b1)
    (D => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b0 && CIX == 1'b1)
    (D => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b1 && CIX == 1'b0)
    (D => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b1 && CIX == 1'b0)
    (D => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b0 && CIX == 1'b1)
    (D => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b0 && CIX == 1'b1)
    (D => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b1 && CIX == 1'b1)
    (D => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b1 && CIX == 1'b1)
    (D => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b0 && CIX == 1'b0)
    (D => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b0 && CIX == 1'b0)
    (D => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DCAP;
    // No function
endmodule
`endcelldefine

`celldefine
module DCAP16;
    // No function
endmodule
`endcelldefine

`celldefine
module DCAP32;
    // No function
endmodule
`endcelldefine

`celldefine
module DCAP4;
    // No function
endmodule
`endcelldefine

`celldefine
module DCAP64;
    // No function
endmodule
`endcelldefine

`celldefine
module DCAP8;
    // No function
endmodule
`endcelldefine

`celldefine
module DEL0 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DEL005 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DEL01 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DEL015 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DEL02 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DEL1 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DEL2 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DEL3 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DEL4 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DFCND1 (D, CP, CDN, Q, QN);
    input D, CP, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, CP_d;
        pullup (SDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCP, CP);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  buf  (CP_check, CDN_i);
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFCND2 (D, CP, CDN, Q, QN);
    input D, CP, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, CP_d;
        pullup (SDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCP, CP);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  buf  (CP_check, CDN_i);
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFCND4 (D, CP, CDN, Q, QN);
    input D, CP, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, CP_d;
        pullup (SDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCP, CP);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  buf  (CP_check, CDN_i);
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFCNQD1 (D, CP, CDN, Q);
    input D, CP, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, CP_d;
        pullup (SDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCP, CP);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  buf  (CP_check, CDN_i);
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFCNQD2 (D, CP, CDN, Q);
    input D, CP, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, CP_d;
        pullup (SDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCP, CP);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  buf  (CP_check, CDN_i);
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFCNQD4 (D, CP, CDN, Q);
    input D, CP, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, CP_d;
        pullup (SDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCP, CP);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  buf  (CP_check, CDN_i);
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFCSND1 (D, CP, CDN, SDN, Q, QN);
    input D, CP, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CP_d;
        tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SDN_SDFCHK, CP_D_SDN, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SDFCHK, CP_nD_SDN, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SDFCHK, nCP_D_SDN, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SDFCHK, nCP_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_CP_D_SDFCHK, CDN_CP_D, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SDFCHK, CDN_CP_nD, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SDFCHK, CDN_nCP_D, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SDFCHK, CDN_nCP_nD, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCP, CP);
    and (CP_D_SDN, CP, D, SDN);
    and (CP_nD_SDN, CP, nD, SDN);
    and (nCP_D_SDN, nCP, D, SDN);
    and (nCP_nD_SDN, nCP, nD, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_CP_D, CDN, CP, D);
    and (CDN_CP_nD, CDN, CP, nD);
    and (CDN_nCP_D, CDN, nCP, D);
    and (CDN_nCP_nD, CDN, nCP, nD);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  and  (CP_check, CDN_i, SDN_i);
  and  (D_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (posedge CP &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (posedge CP &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFCSND2 (D, CP, CDN, SDN, Q, QN);
    input D, CP, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CP_d;
        tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SDN_SDFCHK, CP_D_SDN, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SDFCHK, CP_nD_SDN, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SDFCHK, nCP_D_SDN, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SDFCHK, nCP_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_CP_D_SDFCHK, CDN_CP_D, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SDFCHK, CDN_CP_nD, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SDFCHK, CDN_nCP_D, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SDFCHK, CDN_nCP_nD, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCP, CP);
    and (CP_D_SDN, CP, D, SDN);
    and (CP_nD_SDN, CP, nD, SDN);
    and (nCP_D_SDN, nCP, D, SDN);
    and (nCP_nD_SDN, nCP, nD, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_CP_D, CDN, CP, D);
    and (CDN_CP_nD, CDN, CP, nD);
    and (CDN_nCP_D, CDN, nCP, D);
    and (CDN_nCP_nD, CDN, nCP, nD);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  and  (CP_check, CDN_i, SDN_i);
  and  (D_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (posedge CP &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (posedge CP &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFCSND4 (D, CP, CDN, SDN, Q, QN);
    input D, CP, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CP_d;
        tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SDN_SDFCHK, CP_D_SDN, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SDFCHK, CP_nD_SDN, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SDFCHK, nCP_D_SDN, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SDFCHK, nCP_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_CP_D_SDFCHK, CDN_CP_D, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SDFCHK, CDN_CP_nD, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SDFCHK, CDN_nCP_D, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SDFCHK, CDN_nCP_nD, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCP, CP);
    and (CP_D_SDN, CP, D, SDN);
    and (CP_nD_SDN, CP, nD, SDN);
    and (nCP_D_SDN, nCP, D, SDN);
    and (nCP_nD_SDN, nCP, nD, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_CP_D, CDN, CP, D);
    and (CDN_CP_nD, CDN, CP, nD);
    and (CDN_nCP_D, CDN, nCP, D);
    and (CDN_nCP_nD, CDN, nCP, nD);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  and  (CP_check, CDN_i, SDN_i);
  and  (D_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (posedge CP &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (posedge CP &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFCSNQD1 (D, CP, CDN, SDN, Q);
    input D, CP, CDN, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CP_d;
        tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SDN_SDFCHK, CP_D_SDN, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SDFCHK, CP_nD_SDN, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SDFCHK, nCP_D_SDN, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SDFCHK, nCP_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_CP_D_SDFCHK, CDN_CP_D, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SDFCHK, CDN_CP_nD, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SDFCHK, CDN_nCP_D, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SDFCHK, CDN_nCP_nD, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCP, CP);
    and (CP_D_SDN, CP, D, SDN);
    and (CP_nD_SDN, CP, nD, SDN);
    and (nCP_D_SDN, nCP, D, SDN);
    and (nCP_nD_SDN, nCP, nD, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_CP_D, CDN, CP, D);
    and (CDN_CP_nD, CDN, CP, nD);
    and (CDN_nCP_D, CDN, nCP, D);
    and (CDN_nCP_nD, CDN, nCP, nD);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  and  (CP_check, CDN_i, SDN_i);
  and  (D_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (posedge CP &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (posedge CP &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFCSNQD2 (D, CP, CDN, SDN, Q);
    input D, CP, CDN, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CP_d;
        tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SDN_SDFCHK, CP_D_SDN, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SDFCHK, CP_nD_SDN, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SDFCHK, nCP_D_SDN, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SDFCHK, nCP_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_CP_D_SDFCHK, CDN_CP_D, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SDFCHK, CDN_CP_nD, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SDFCHK, CDN_nCP_D, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SDFCHK, CDN_nCP_nD, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCP, CP);
    and (CP_D_SDN, CP, D, SDN);
    and (CP_nD_SDN, CP, nD, SDN);
    and (nCP_D_SDN, nCP, D, SDN);
    and (nCP_nD_SDN, nCP, nD, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_CP_D, CDN, CP, D);
    and (CDN_CP_nD, CDN, CP, nD);
    and (CDN_nCP_D, CDN, nCP, D);
    and (CDN_nCP_nD, CDN, nCP, nD);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  and  (CP_check, CDN_i, SDN_i);
  and  (D_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (posedge CP &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (posedge CP &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFCSNQD4 (D, CP, CDN, SDN, Q);
    input D, CP, CDN, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CP_d;
        tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SDN_SDFCHK, CP_D_SDN, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SDFCHK, CP_nD_SDN, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SDFCHK, nCP_D_SDN, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SDFCHK, nCP_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_CP_D_SDFCHK, CDN_CP_D, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SDFCHK, CDN_CP_nD, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SDFCHK, CDN_nCP_D, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SDFCHK, CDN_nCP_nD, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCP, CP);
    and (CP_D_SDN, CP, D, SDN);
    and (CP_nD_SDN, CP, nD, SDN);
    and (nCP_D_SDN, nCP, D, SDN);
    and (nCP_nD_SDN, nCP, nD, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_CP_D, CDN, CP, D);
    and (CDN_CP_nD, CDN, CP, nD);
    and (CDN_nCP_D, CDN, nCP, D);
    and (CDN_nCP_nD, CDN, nCP, nD);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  and  (CP_check, CDN_i, SDN_i);
  and  (D_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (posedge CP &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (posedge CP &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFD1 (D, CP, Q, QN);
    input D, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
  `endif

    not (nD, D);

  // Timing logics defined for default constraint check
  pullup  (CP_check);
  pullup  (D_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:D)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    $width (posedge CP &&& D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFD2 (D, CP, Q, QN);
    input D, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
  `endif

    not (nD, D);

  // Timing logics defined for default constraint check
  pullup  (CP_check);
  pullup  (D_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:D)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    $width (posedge CP &&& D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFD4 (D, CP, Q, QN);
    input D, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
  `endif

    not (nD, D);

  // Timing logics defined for default constraint check
  pullup  (CP_check);
  pullup  (D_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:D)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    $width (posedge CP &&& D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKCND1 (D, CP, CN, Q, QN);
    input D, CP, CN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        and (D_i, CN_d, D_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        and (D_i, CN, D);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (CN_SDFCHK, CN, 1'b1);
    tsmc_xbuf (CN_D_SDFCHK, CN_D, 1'b1);
    tsmc_xbuf (CN_nD_SDFCHK, CN_nD, 1'b1);
    tsmc_xbuf (nCN_D_SDFCHK, nCN_D, 1'b1);
    tsmc_xbuf (nCN_nD_SDFCHK, nCN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCN, CN);
    and (CN_D, CN, D);
    and (CN_nD, CN, nD);
    and (nCN_D, nCN, D);
    and (nCN_nD, nCN, nD);

  // Timing logics defined for default constraint check
  `ifdef NTC
    buf  (D_check, CN_d);
  `else
    buf  (D_check, CN);
  `endif
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((CN && D)))) = (0, 0);
    (posedge CP => (QN-:((CN && D)))) = (0, 0);
    $width (posedge CP &&& CN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP &&& D_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SDFCHK, negedge D , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKCND2 (D, CP, CN, Q, QN);
    input D, CP, CN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        and (D_i, CN_d, D_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        and (D_i, CN, D);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (CN_SDFCHK, CN, 1'b1);
    tsmc_xbuf (CN_D_SDFCHK, CN_D, 1'b1);
    tsmc_xbuf (CN_nD_SDFCHK, CN_nD, 1'b1);
    tsmc_xbuf (nCN_D_SDFCHK, nCN_D, 1'b1);
    tsmc_xbuf (nCN_nD_SDFCHK, nCN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCN, CN);
    and (CN_D, CN, D);
    and (CN_nD, CN, nD);
    and (nCN_D, nCN, D);
    and (nCN_nD, nCN, nD);

  // Timing logics defined for default constraint check
  `ifdef NTC
    buf  (D_check, CN_d);
  `else
    buf  (D_check, CN);
  `endif
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((CN && D)))) = (0, 0);
    (posedge CP => (QN-:((CN && D)))) = (0, 0);
    $width (posedge CP &&& CN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP &&& D_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SDFCHK, negedge D , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKCND4 (D, CP, CN, Q, QN);
    input D, CP, CN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        and (D_i, CN_d, D_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        and (D_i, CN, D);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (CN_SDFCHK, CN, 1'b1);
    tsmc_xbuf (CN_D_SDFCHK, CN_D, 1'b1);
    tsmc_xbuf (CN_nD_SDFCHK, CN_nD, 1'b1);
    tsmc_xbuf (nCN_D_SDFCHK, nCN_D, 1'b1);
    tsmc_xbuf (nCN_nD_SDFCHK, nCN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCN, CN);
    and (CN_D, CN, D);
    and (CN_nD, CN, nD);
    and (nCN_D, nCN, D);
    and (nCN_nD, nCN, nD);

  // Timing logics defined for default constraint check
  `ifdef NTC
    buf  (D_check, CN_d);
  `else
    buf  (D_check, CN);
  `endif
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((CN && D)))) = (0, 0);
    (posedge CP => (QN-:((CN && D)))) = (0, 0);
    $width (posedge CP &&& CN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP &&& D_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SDFCHK, negedge D , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKCNQD1 (D, CP, CN, Q);
    input D, CP, CN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        and (D_i, CN_d, D_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        and (D_i, CN, D);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (CN_SDFCHK, CN, 1'b1);
    tsmc_xbuf (CN_D_SDFCHK, CN_D, 1'b1);
    tsmc_xbuf (CN_nD_SDFCHK, CN_nD, 1'b1);
    tsmc_xbuf (nCN_D_SDFCHK, nCN_D, 1'b1);
    tsmc_xbuf (nCN_nD_SDFCHK, nCN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCN, CN);
    and (CN_D, CN, D);
    and (CN_nD, CN, nD);
    and (nCN_D, nCN, D);
    and (nCN_nD, nCN, nD);

  // Timing logics defined for default constraint check
  `ifdef NTC
    buf  (D_check, CN_d);
  `else
    buf  (D_check, CN);
  `endif
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((CN && D)))) = (0, 0);
    $width (posedge CP &&& CN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP &&& D_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SDFCHK, negedge D , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKCNQD2 (D, CP, CN, Q);
    input D, CP, CN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        and (D_i, CN_d, D_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        and (D_i, CN, D);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (CN_SDFCHK, CN, 1'b1);
    tsmc_xbuf (CN_D_SDFCHK, CN_D, 1'b1);
    tsmc_xbuf (CN_nD_SDFCHK, CN_nD, 1'b1);
    tsmc_xbuf (nCN_D_SDFCHK, nCN_D, 1'b1);
    tsmc_xbuf (nCN_nD_SDFCHK, nCN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCN, CN);
    and (CN_D, CN, D);
    and (CN_nD, CN, nD);
    and (nCN_D, nCN, D);
    and (nCN_nD, nCN, nD);

  // Timing logics defined for default constraint check
  `ifdef NTC
    buf  (D_check, CN_d);
  `else
    buf  (D_check, CN);
  `endif
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((CN && D)))) = (0, 0);
    $width (posedge CP &&& CN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP &&& D_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SDFCHK, negedge D , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKCNQD4 (D, CP, CN, Q);
    input D, CP, CN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        and (D_i, CN_d, D_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        and (D_i, CN, D);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (CN_SDFCHK, CN, 1'b1);
    tsmc_xbuf (CN_D_SDFCHK, CN_D, 1'b1);
    tsmc_xbuf (CN_nD_SDFCHK, CN_nD, 1'b1);
    tsmc_xbuf (nCN_D_SDFCHK, nCN_D, 1'b1);
    tsmc_xbuf (nCN_nD_SDFCHK, nCN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCN, CN);
    and (CN_D, CN, D);
    and (CN_nD, CN, nD);
    and (nCN_D, nCN, D);
    and (nCN_nD, nCN, nD);

  // Timing logics defined for default constraint check
  `ifdef NTC
    buf  (D_check, CN_d);
  `else
    buf  (D_check, CN);
  `endif
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((CN && D)))) = (0, 0);
    $width (posedge CP &&& CN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP &&& D_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SDFCHK, negedge D , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKCSND1 (D, CP, CN, SN, Q, QN);
    input D, CP, CN, SN;
    output Q, QN;
    reg notifier;
    reg flag;
    `ifdef NTC
        wire D_d, CP_d, CN_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (DS, S, D_d);
        and (D_i, CN_d, DS);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (DS, S, D);
        and (D_i, CN, DS);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 
    buf (CN_i, CN);
    buf (SN_i, SN);
    always @(CN_i or SN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CN_i===1'b0)&&(SN_i===1'b0));
            if (flag == 1) begin 
                if (CN_i!==1'b0) begin
                    $display("%m > CN is released at time %.2fns.", $realtime);
                end 
                if (SN_i!==1'b0) begin
                    $display("%m > SN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CN and SN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SN_SDFCHK, CN_D_SN, 1'b1);
    tsmc_xbuf (CN_D_nSN_SDFCHK, CN_D_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSN_SDFCHK, CN_nD_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SN_SDFCHK, CN_nD_SN, 1'b1);
    tsmc_xbuf (nCN_D_SN_SDFCHK, nCN_D_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SN_SDFCHK, nCN_nD_SN, 1'b1);
    tsmc_xbuf (D_SN_SDFCHK, D_SN, 1'b1);
    tsmc_xbuf (CN_SN_SDFCHK, CN_SN, 1'b1);
    tsmc_xbuf (CN_nD_SDFCHK, CN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCN, CN);
    not (nSN, SN);
    and (CN_D_SN, CN, D, SN);
    and (CN_D_nSN, CN, D, nSN);
    and (CN_nD_nSN, CN, nD, nSN);
    and (CN_nD_SN, CN, nD, SN);
    and (nCN_D_SN, nCN, D, SN);
    and (nCN_nD_SN, nCN, nD, SN);
    and (D_SN, D, SN);
    and (CN_SN, CN, SN);
    and (CN_nD, CN, nD);

  // Timing logics defined for default constraint check
  `ifdef NTC
    buf  (SN_check, CN_d);
    and  (D_check, SN_d, CN_d);
  `else
    buf  (SN_check, CN);
    and  (D_check, SN, CN);
  `endif
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((CN && D) || (CN && !(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((CN && D) || (CN && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& CN_D_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& D_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKCSND2 (D, CP, CN, SN, Q, QN);
    input D, CP, CN, SN;
    output Q, QN;
    reg notifier;
    reg flag;
    `ifdef NTC
        wire D_d, CP_d, CN_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (DS, S, D_d);
        and (D_i, CN_d, DS);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (DS, S, D);
        and (D_i, CN, DS);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 
    buf (CN_i, CN);
    buf (SN_i, SN);
    always @(CN_i or SN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CN_i===1'b0)&&(SN_i===1'b0));
            if (flag == 1) begin 
                if (CN_i!==1'b0) begin
                    $display("%m > CN is released at time %.2fns.", $realtime);
                end 
                if (SN_i!==1'b0) begin
                    $display("%m > SN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CN and SN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SN_SDFCHK, CN_D_SN, 1'b1);
    tsmc_xbuf (CN_D_nSN_SDFCHK, CN_D_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSN_SDFCHK, CN_nD_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SN_SDFCHK, CN_nD_SN, 1'b1);
    tsmc_xbuf (nCN_D_SN_SDFCHK, nCN_D_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SN_SDFCHK, nCN_nD_SN, 1'b1);
    tsmc_xbuf (D_SN_SDFCHK, D_SN, 1'b1);
    tsmc_xbuf (CN_SN_SDFCHK, CN_SN, 1'b1);
    tsmc_xbuf (CN_nD_SDFCHK, CN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCN, CN);
    not (nSN, SN);
    and (CN_D_SN, CN, D, SN);
    and (CN_D_nSN, CN, D, nSN);
    and (CN_nD_nSN, CN, nD, nSN);
    and (CN_nD_SN, CN, nD, SN);
    and (nCN_D_SN, nCN, D, SN);
    and (nCN_nD_SN, nCN, nD, SN);
    and (D_SN, D, SN);
    and (CN_SN, CN, SN);
    and (CN_nD, CN, nD);

  // Timing logics defined for default constraint check
  `ifdef NTC
    buf  (SN_check, CN_d);
    and  (D_check, SN_d, CN_d);
  `else
    buf  (SN_check, CN);
    and  (D_check, SN, CN);
  `endif
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((CN && D) || (CN && !(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((CN && D) || (CN && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& CN_D_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& D_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKCSND4 (D, CP, CN, SN, Q, QN);
    input D, CP, CN, SN;
    output Q, QN;
    reg notifier;
    reg flag;
    `ifdef NTC
        wire D_d, CP_d, CN_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (DS, S, D_d);
        and (D_i, CN_d, DS);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (DS, S, D);
        and (D_i, CN, DS);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 
    buf (CN_i, CN);
    buf (SN_i, SN);
    always @(CN_i or SN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CN_i===1'b0)&&(SN_i===1'b0));
            if (flag == 1) begin 
                if (CN_i!==1'b0) begin
                    $display("%m > CN is released at time %.2fns.", $realtime);
                end 
                if (SN_i!==1'b0) begin
                    $display("%m > SN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CN and SN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SN_SDFCHK, CN_D_SN, 1'b1);
    tsmc_xbuf (CN_D_nSN_SDFCHK, CN_D_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSN_SDFCHK, CN_nD_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SN_SDFCHK, CN_nD_SN, 1'b1);
    tsmc_xbuf (nCN_D_SN_SDFCHK, nCN_D_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SN_SDFCHK, nCN_nD_SN, 1'b1);
    tsmc_xbuf (D_SN_SDFCHK, D_SN, 1'b1);
    tsmc_xbuf (CN_SN_SDFCHK, CN_SN, 1'b1);
    tsmc_xbuf (CN_nD_SDFCHK, CN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCN, CN);
    not (nSN, SN);
    and (CN_D_SN, CN, D, SN);
    and (CN_D_nSN, CN, D, nSN);
    and (CN_nD_nSN, CN, nD, nSN);
    and (CN_nD_SN, CN, nD, SN);
    and (nCN_D_SN, nCN, D, SN);
    and (nCN_nD_SN, nCN, nD, SN);
    and (D_SN, D, SN);
    and (CN_SN, CN, SN);
    and (CN_nD, CN, nD);

  // Timing logics defined for default constraint check
  `ifdef NTC
    buf  (SN_check, CN_d);
    and  (D_check, SN_d, CN_d);
  `else
    buf  (SN_check, CN);
    and  (D_check, SN, CN);
  `endif
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((CN && D) || (CN && !(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((CN && D) || (CN && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& CN_D_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& D_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKSND1 (D, CP, SN, Q, QN);
    input D, CP, SN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (D_i, S, D_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (D_i, S, D);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SN_SDFCHK, SN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SN_SDFCHK, D_SN, 1'b1);
    tsmc_xbuf (D_nSN_SDFCHK, D_nSN, 1'b1);
    tsmc_xbuf (nD_nSN_SDFCHK, nD_nSN, 1'b1);
    tsmc_xbuf (nD_SN_SDFCHK, nD_SN, 1'b1);
  `endif

    not (nD, D);
    not (nSN, SN);
    and (D_SN, D, SN);
    and (D_nSN, D, nSN);
    and (nD_nSN, nD, nSN);
    and (nD_SN, nD, SN);

  // Timing logics defined for default constraint check
  `ifdef NTC
    buf  (D_check, SN_d);
  `else
    buf  (D_check, SN);
  `endif
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((D) || (!(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((D) || (!(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& D_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKSND2 (D, CP, SN, Q, QN);
    input D, CP, SN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (D_i, S, D_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (D_i, S, D);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SN_SDFCHK, SN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SN_SDFCHK, D_SN, 1'b1);
    tsmc_xbuf (D_nSN_SDFCHK, D_nSN, 1'b1);
    tsmc_xbuf (nD_nSN_SDFCHK, nD_nSN, 1'b1);
    tsmc_xbuf (nD_SN_SDFCHK, nD_SN, 1'b1);
  `endif

    not (nD, D);
    not (nSN, SN);
    and (D_SN, D, SN);
    and (D_nSN, D, nSN);
    and (nD_nSN, nD, nSN);
    and (nD_SN, nD, SN);

  // Timing logics defined for default constraint check
  `ifdef NTC
    buf  (D_check, SN_d);
  `else
    buf  (D_check, SN);
  `endif
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((D) || (!(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((D) || (!(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& D_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKSND4 (D, CP, SN, Q, QN);
    input D, CP, SN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (D_i, S, D_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (D_i, S, D);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SN_SDFCHK, SN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SN_SDFCHK, D_SN, 1'b1);
    tsmc_xbuf (D_nSN_SDFCHK, D_nSN, 1'b1);
    tsmc_xbuf (nD_nSN_SDFCHK, nD_nSN, 1'b1);
    tsmc_xbuf (nD_SN_SDFCHK, nD_SN, 1'b1);
  `endif

    not (nD, D);
    not (nSN, SN);
    and (D_SN, D, SN);
    and (D_nSN, D, nSN);
    and (nD_nSN, nD, nSN);
    and (nD_SN, nD, SN);

  // Timing logics defined for default constraint check
  `ifdef NTC
    buf  (D_check, SN_d);
  `else
    buf  (D_check, SN);
  `endif
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((D) || (!(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((D) || (!(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& D_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFNCND1 (D, CPN, CDN, Q, QN);
    input D, CPN, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, CPN_d;
        pullup (SDN);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_d, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        not (CP, CPN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (CPN_D_SDFCHK, CPN_D, 1'b1);
    tsmc_xbuf (CPN_nD_SDFCHK, CPN_nD, 1'b1);
    tsmc_xbuf (nCPN_D_SDFCHK, nCPN_D, 1'b1);
    tsmc_xbuf (nCPN_nD_SDFCHK, nCPN_nD, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCPN, CPN);
    and (CPN_D, CPN, D);
    and (CPN_nD, CPN, nD);
    and (nCPN_D, nCPN, D);
    and (nCPN_nD, nCPN, nD);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  buf  (CPN_check, CDN_i);
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CPN == 1'b1 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:D)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    $width (negedge CDN &&& CPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, negedge CPN &&& D_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, negedge CPN &&& D_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, negedge CPN &&& D_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFNCND2 (D, CPN, CDN, Q, QN);
    input D, CPN, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, CPN_d;
        pullup (SDN);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_d, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        not (CP, CPN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (CPN_D_SDFCHK, CPN_D, 1'b1);
    tsmc_xbuf (CPN_nD_SDFCHK, CPN_nD, 1'b1);
    tsmc_xbuf (nCPN_D_SDFCHK, nCPN_D, 1'b1);
    tsmc_xbuf (nCPN_nD_SDFCHK, nCPN_nD, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCPN, CPN);
    and (CPN_D, CPN, D);
    and (CPN_nD, CPN, nD);
    and (nCPN_D, nCPN, D);
    and (nCPN_nD, nCPN, nD);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  buf  (CPN_check, CDN_i);
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CPN == 1'b1 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:D)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    $width (negedge CDN &&& CPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, negedge CPN &&& D_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, negedge CPN &&& D_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, negedge CPN &&& D_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFNCND4 (D, CPN, CDN, Q, QN);
    input D, CPN, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, CPN_d;
        pullup (SDN);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_d, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        not (CP, CPN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (CPN_D_SDFCHK, CPN_D, 1'b1);
    tsmc_xbuf (CPN_nD_SDFCHK, CPN_nD, 1'b1);
    tsmc_xbuf (nCPN_D_SDFCHK, nCPN_D, 1'b1);
    tsmc_xbuf (nCPN_nD_SDFCHK, nCPN_nD, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCPN, CPN);
    and (CPN_D, CPN, D);
    and (CPN_nD, CPN, nD);
    and (nCPN_D, nCPN, D);
    and (nCPN_nD, nCPN, nD);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  buf  (CPN_check, CDN_i);
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CPN == 1'b1 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:D)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    $width (negedge CDN &&& CPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, negedge CPN &&& D_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, negedge CPN &&& D_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, negedge CPN &&& D_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFNCSND1 (D, CPN, CDN, SDN, Q, QN);
    input D, CPN, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CPN_d;
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_d, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        not (CP, CPN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_D_SDN_SDFCHK, CPN_D_SDN, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_SDFCHK, CPN_nD_SDN, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_SDFCHK, nCPN_D_SDN, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_SDFCHK, nCPN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_CPN_D_SDFCHK, CDN_CPN_D, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_SDFCHK, CDN_CPN_nD, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_SDFCHK, CDN_nCPN_D, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_SDFCHK, CDN_nCPN_nD, 1'b1);
    tsmc_xbuf (CPN_D_SDFCHK, CPN_D, 1'b1);
    tsmc_xbuf (CPN_nD_SDFCHK, CPN_nD, 1'b1);
    tsmc_xbuf (nCPN_D_SDFCHK, nCPN_D, 1'b1);
    tsmc_xbuf (nCPN_nD_SDFCHK, nCPN_nD, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCPN, CPN);
    and (CPN_D_SDN, CPN, D, SDN);
    and (CPN_nD_SDN, CPN, nD, SDN);
    and (nCPN_D_SDN, nCPN, D, SDN);
    and (nCPN_nD_SDN, nCPN, nD, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_CPN_D, CDN, CPN, D);
    and (CDN_CPN_nD, CDN, CPN, nD);
    and (CDN_nCPN_D, CDN, nCPN, D);
    and (CDN_nCPN_nD, CDN, nCPN, nD);
    and (CPN_D, CPN, D);
    and (CPN_nD, CPN, nD);
    and (nCPN_D, nCPN, D);
    and (nCPN_nD, nCPN, nD);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  and  (CPN_check, CDN_i, SDN_i);
  and  (D_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge CDN &&& CPN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CPN_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (posedge CDN &&& CPN_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, negedge CPN &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, negedge CPN &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (posedge SDN &&& CPN_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (posedge CDN &&& CPN_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge CPN &&& D_SDN_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge CPN &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CPN_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge CPN &&& D_SDN_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge CPN &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFNCSND2 (D, CPN, CDN, SDN, Q, QN);
    input D, CPN, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CPN_d;
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_d, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        not (CP, CPN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_D_SDN_SDFCHK, CPN_D_SDN, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_SDFCHK, CPN_nD_SDN, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_SDFCHK, nCPN_D_SDN, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_SDFCHK, nCPN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_CPN_D_SDFCHK, CDN_CPN_D, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_SDFCHK, CDN_CPN_nD, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_SDFCHK, CDN_nCPN_D, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_SDFCHK, CDN_nCPN_nD, 1'b1);
    tsmc_xbuf (CPN_D_SDFCHK, CPN_D, 1'b1);
    tsmc_xbuf (CPN_nD_SDFCHK, CPN_nD, 1'b1);
    tsmc_xbuf (nCPN_D_SDFCHK, nCPN_D, 1'b1);
    tsmc_xbuf (nCPN_nD_SDFCHK, nCPN_nD, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCPN, CPN);
    and (CPN_D_SDN, CPN, D, SDN);
    and (CPN_nD_SDN, CPN, nD, SDN);
    and (nCPN_D_SDN, nCPN, D, SDN);
    and (nCPN_nD_SDN, nCPN, nD, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_CPN_D, CDN, CPN, D);
    and (CDN_CPN_nD, CDN, CPN, nD);
    and (CDN_nCPN_D, CDN, nCPN, D);
    and (CDN_nCPN_nD, CDN, nCPN, nD);
    and (CPN_D, CPN, D);
    and (CPN_nD, CPN, nD);
    and (nCPN_D, nCPN, D);
    and (nCPN_nD, nCPN, nD);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  and  (CPN_check, CDN_i, SDN_i);
  and  (D_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge CDN &&& CPN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CPN_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (posedge CDN &&& CPN_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, negedge CPN &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, negedge CPN &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (posedge SDN &&& CPN_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (posedge CDN &&& CPN_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge CPN &&& D_SDN_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge CPN &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CPN_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge CPN &&& D_SDN_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge CPN &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFNCSND4 (D, CPN, CDN, SDN, Q, QN);
    input D, CPN, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CPN_d;
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_d, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        not (CP, CPN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_D_SDN_SDFCHK, CPN_D_SDN, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_SDFCHK, CPN_nD_SDN, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_SDFCHK, nCPN_D_SDN, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_SDFCHK, nCPN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_CPN_D_SDFCHK, CDN_CPN_D, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_SDFCHK, CDN_CPN_nD, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_SDFCHK, CDN_nCPN_D, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_SDFCHK, CDN_nCPN_nD, 1'b1);
    tsmc_xbuf (CPN_D_SDFCHK, CPN_D, 1'b1);
    tsmc_xbuf (CPN_nD_SDFCHK, CPN_nD, 1'b1);
    tsmc_xbuf (nCPN_D_SDFCHK, nCPN_D, 1'b1);
    tsmc_xbuf (nCPN_nD_SDFCHK, nCPN_nD, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCPN, CPN);
    and (CPN_D_SDN, CPN, D, SDN);
    and (CPN_nD_SDN, CPN, nD, SDN);
    and (nCPN_D_SDN, nCPN, D, SDN);
    and (nCPN_nD_SDN, nCPN, nD, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_CPN_D, CDN, CPN, D);
    and (CDN_CPN_nD, CDN, CPN, nD);
    and (CDN_nCPN_D, CDN, nCPN, D);
    and (CDN_nCPN_nD, CDN, nCPN, nD);
    and (CPN_D, CPN, D);
    and (CPN_nD, CPN, nD);
    and (nCPN_D, nCPN, D);
    and (nCPN_nD, nCPN, nD);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  and  (CPN_check, CDN_i, SDN_i);
  and  (D_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge CDN &&& CPN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CPN_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (posedge CDN &&& CPN_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, negedge CPN &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, negedge CPN &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (posedge SDN &&& CPN_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (posedge CDN &&& CPN_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge CPN &&& D_SDN_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge CPN &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CPN_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge CPN &&& D_SDN_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge CPN &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFND1 (D, CPN, Q, QN);
    input D, CPN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, CPN_d;
        pullup (CDN);
        pullup (SDN);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_d, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (CP, CPN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
  `endif

    not (nD, D);

  // Timing logics defined for default constraint check
  pullup  (CPN_check);
  pullup  (D_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CPN => (Q+:D)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    $width (posedge CPN &&& D_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
  `else
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFND2 (D, CPN, Q, QN);
    input D, CPN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, CPN_d;
        pullup (CDN);
        pullup (SDN);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_d, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (CP, CPN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
  `endif

    not (nD, D);

  // Timing logics defined for default constraint check
  pullup  (CPN_check);
  pullup  (D_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CPN => (Q+:D)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    $width (posedge CPN &&& D_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
  `else
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFND4 (D, CPN, Q, QN);
    input D, CPN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, CPN_d;
        pullup (CDN);
        pullup (SDN);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_d, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (CP, CPN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
  `endif

    not (nD, D);

  // Timing logics defined for default constraint check
  pullup  (CPN_check);
  pullup  (D_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CPN => (Q+:D)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    $width (posedge CPN &&& D_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
  `else
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFNSND1 (D, CPN, SDN, Q, QN);
    input D, CPN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CPN_d;
        pullup (CDN);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_d, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        not (CP, CPN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (CPN_D_SDFCHK, CPN_D, 1'b1);
    tsmc_xbuf (CPN_nD_SDFCHK, CPN_nD, 1'b1);
    tsmc_xbuf (nCPN_D_SDFCHK, nCPN_D, 1'b1);
    tsmc_xbuf (nCPN_nD_SDFCHK, nCPN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCPN, CPN);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (CPN_D, CPN, D);
    and (CPN_nD, CPN, nD);
    and (nCPN_D, nCPN, D);
    and (nCPN_nD, nCPN, nD);

  // Timing logics defined for default constraint check
  buf  (CPN_check, SDN_i);
  buf  (D_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CPN => (Q+:D)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CPN &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, negedge CPN &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, negedge CPN &&& nD_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, negedge CPN &&& nD_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFNSND2 (D, CPN, SDN, Q, QN);
    input D, CPN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CPN_d;
        pullup (CDN);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_d, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        not (CP, CPN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (CPN_D_SDFCHK, CPN_D, 1'b1);
    tsmc_xbuf (CPN_nD_SDFCHK, CPN_nD, 1'b1);
    tsmc_xbuf (nCPN_D_SDFCHK, nCPN_D, 1'b1);
    tsmc_xbuf (nCPN_nD_SDFCHK, nCPN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCPN, CPN);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (CPN_D, CPN, D);
    and (CPN_nD, CPN, nD);
    and (nCPN_D, nCPN, D);
    and (nCPN_nD, nCPN, nD);

  // Timing logics defined for default constraint check
  buf  (CPN_check, SDN_i);
  buf  (D_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CPN => (Q+:D)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CPN &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, negedge CPN &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, negedge CPN &&& nD_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, negedge CPN &&& nD_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFNSND4 (D, CPN, SDN, Q, QN);
    input D, CPN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CPN_d;
        pullup (CDN);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_d, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        not (CP, CPN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (CPN_D_SDFCHK, CPN_D, 1'b1);
    tsmc_xbuf (CPN_nD_SDFCHK, CPN_nD, 1'b1);
    tsmc_xbuf (nCPN_D_SDFCHK, nCPN_D, 1'b1);
    tsmc_xbuf (nCPN_nD_SDFCHK, nCPN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCPN, CPN);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (CPN_D, CPN, D);
    and (CPN_nD, CPN, nD);
    and (nCPN_D, nCPN, D);
    and (nCPN_nD, nCPN, nD);

  // Timing logics defined for default constraint check
  buf  (CPN_check, SDN_i);
  buf  (D_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CPN => (Q+:D)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CPN &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, negedge CPN &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, negedge CPN &&& nD_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, negedge CPN &&& nD_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFQD1 (D, CP, Q);
    input D, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
  `endif

    not (nD, D);

  // Timing logics defined for default constraint check
  pullup  (CP_check);
  pullup  (D_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:D)) = (0, 0);
    $width (posedge CP &&& D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFQD2 (D, CP, Q);
    input D, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
  `endif

    not (nD, D);

  // Timing logics defined for default constraint check
  pullup  (CP_check);
  pullup  (D_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:D)) = (0, 0);
    $width (posedge CP &&& D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFQD4 (D, CP, Q);
    input D, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
  `endif

    not (nD, D);

  // Timing logics defined for default constraint check
  pullup  (CP_check);
  pullup  (D_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:D)) = (0, 0);
    $width (posedge CP &&& D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFSND1 (D, CP, SDN, Q, QN);
    input D, CP, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CP_d;
        pullup (CDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCP, CP);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);

  // Timing logics defined for default constraint check
  buf  (CP_check, SDN_i);
  buf  (D_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:D)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0, notifier);
      $hold (posedge CP &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0, notifier);
    $hold (posedge CP &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFSND2 (D, CP, SDN, Q, QN);
    input D, CP, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CP_d;
        pullup (CDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCP, CP);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);

  // Timing logics defined for default constraint check
  buf  (CP_check, SDN_i);
  buf  (D_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:D)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0, notifier);
      $hold (posedge CP &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0, notifier);
    $hold (posedge CP &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFSND4 (D, CP, SDN, Q, QN);
    input D, CP, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CP_d;
        pullup (CDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCP, CP);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);

  // Timing logics defined for default constraint check
  buf  (CP_check, SDN_i);
  buf  (D_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:D)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0, notifier);
      $hold (posedge CP &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0, notifier);
    $hold (posedge CP &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFSNQD1 (D, CP, SDN, Q);
    input D, CP, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CP_d;
        pullup (CDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCP, CP);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);

  // Timing logics defined for default constraint check
  buf  (CP_check, SDN_i);
  buf  (D_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:D)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0, notifier);
      $hold (posedge CP &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0, notifier);
    $hold (posedge CP &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFSNQD2 (D, CP, SDN, Q);
    input D, CP, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CP_d;
        pullup (CDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCP, CP);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);

  // Timing logics defined for default constraint check
  buf  (CP_check, SDN_i);
  buf  (D_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:D)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0, notifier);
      $hold (posedge CP &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0, notifier);
    $hold (posedge CP &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFSNQD4 (D, CP, SDN, Q);
    input D, CP, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CP_d;
        pullup (CDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
  `endif

    not (nD, D);
    not (nCP, CP);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);

  // Timing logics defined for default constraint check
  buf  (CP_check, SDN_i);
  buf  (D_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:D)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0, notifier);
      $hold (posedge CP &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0, notifier);
    $hold (posedge CP &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFXD1 (DA, DB, SA, CP, Q, QN);
    input DA, DB, SA, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire DA_d, DB_d, SA_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB_d, DA_d, SA_d);
        tsmc_dff (Q_buf, D, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB, DA, SA);
        tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (DA_DB_SA_SDFCHK, DA_DB_SA, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SDFCHK, DA_DB_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SDFCHK, DA_nDB_SA, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SDFCHK, nDA_DB_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SDFCHK, DA_nDB_nSA, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SDFCHK, nDA_DB_SA, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SDFCHK, nDA_nDB_SA, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SDFCHK, nDA_nDB_nSA, 1'b1);
    tsmc_xbuf (DB_SA_SDFCHK, DB_SA, 1'b1);
    tsmc_xbuf (nDB_SA_SDFCHK, nDB_SA, 1'b1);
    tsmc_xbuf (DA_nSA_SDFCHK, DA_nSA, 1'b1);
    tsmc_xbuf (nDA_nSA_SDFCHK, nDA_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_SDFCHK, DA_nDB, 1'b1);
    tsmc_xbuf (nDA_DB_SDFCHK, nDA_DB, 1'b1);
  `endif

    not (nDA, DA);
    not (nDB, DB);
    not (nSA, SA);
    and (DA_DB_SA, DA, DB, SA);
    and (DA_DB_nSA, DA, DB, nSA);
    and (DA_nDB_SA, DA, nDB, SA);
    and (nDA_DB_nSA, nDA, DB, nSA);
    and (DA_nDB_nSA, DA, nDB, nSA);
    and (nDA_DB_SA, nDA, DB, SA);
    and (nDA_nDB_SA, nDA, nDB, SA);
    and (nDA_nDB_nSA, nDA, nDB, nSA);
    and (DB_SA, DB, SA);
    and (nDB_SA, nDB, SA);
    and (DA_nSA, DA, nSA);
    and (nDA_nSA, nDA, nSA);
    and (DA_nDB, DA, nDB);
    and (nDA_DB, nDA, DB);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SA_int_not, SA_d);
    buf  (DA_check, SA_d);
  `else
    not  (SA_int_not, SA);
    buf  (DA_check, SA);
  `endif
  buf  (DB_check, SA_int_not);
  pullup  (CP_check);
  pullup  (SA_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((DA && DB) || (DA && !(DB) && SA) || (!(DA) && DB && !(SA))))) = (0, 0);
    (posedge CP => (QN-:((DA && DB) || (DA && !(DB) && SA) || (!(DA) && DB && !(SA))))) = (0, 0);
    $width (posedge CP &&& DA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DB_SA_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
  `else
    $setuphold (posedge CP &&& DB_SA_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, negedge SA , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFXD2 (DA, DB, SA, CP, Q, QN);
    input DA, DB, SA, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire DA_d, DB_d, SA_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB_d, DA_d, SA_d);
        tsmc_dff (Q_buf, D, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB, DA, SA);
        tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (DA_DB_SA_SDFCHK, DA_DB_SA, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SDFCHK, DA_DB_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SDFCHK, DA_nDB_SA, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SDFCHK, nDA_DB_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SDFCHK, DA_nDB_nSA, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SDFCHK, nDA_DB_SA, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SDFCHK, nDA_nDB_SA, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SDFCHK, nDA_nDB_nSA, 1'b1);
    tsmc_xbuf (DB_SA_SDFCHK, DB_SA, 1'b1);
    tsmc_xbuf (nDB_SA_SDFCHK, nDB_SA, 1'b1);
    tsmc_xbuf (DA_nSA_SDFCHK, DA_nSA, 1'b1);
    tsmc_xbuf (nDA_nSA_SDFCHK, nDA_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_SDFCHK, DA_nDB, 1'b1);
    tsmc_xbuf (nDA_DB_SDFCHK, nDA_DB, 1'b1);
  `endif

    not (nDA, DA);
    not (nDB, DB);
    not (nSA, SA);
    and (DA_DB_SA, DA, DB, SA);
    and (DA_DB_nSA, DA, DB, nSA);
    and (DA_nDB_SA, DA, nDB, SA);
    and (nDA_DB_nSA, nDA, DB, nSA);
    and (DA_nDB_nSA, DA, nDB, nSA);
    and (nDA_DB_SA, nDA, DB, SA);
    and (nDA_nDB_SA, nDA, nDB, SA);
    and (nDA_nDB_nSA, nDA, nDB, nSA);
    and (DB_SA, DB, SA);
    and (nDB_SA, nDB, SA);
    and (DA_nSA, DA, nSA);
    and (nDA_nSA, nDA, nSA);
    and (DA_nDB, DA, nDB);
    and (nDA_DB, nDA, DB);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SA_int_not, SA_d);
    buf  (DA_check, SA_d);
  `else
    not  (SA_int_not, SA);
    buf  (DA_check, SA);
  `endif
  buf  (DB_check, SA_int_not);
  pullup  (CP_check);
  pullup  (SA_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((DA && DB) || (DA && !(DB) && SA) || (!(DA) && DB && !(SA))))) = (0, 0);
    (posedge CP => (QN-:((DA && DB) || (DA && !(DB) && SA) || (!(DA) && DB && !(SA))))) = (0, 0);
    $width (posedge CP &&& DA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DB_SA_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
  `else
    $setuphold (posedge CP &&& DB_SA_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, negedge SA , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFXD4 (DA, DB, SA, CP, Q, QN);
    input DA, DB, SA, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire DA_d, DB_d, SA_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB_d, DA_d, SA_d);
        tsmc_dff (Q_buf, D, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB, DA, SA);
        tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (DA_DB_SA_SDFCHK, DA_DB_SA, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SDFCHK, DA_DB_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SDFCHK, DA_nDB_SA, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SDFCHK, nDA_DB_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SDFCHK, DA_nDB_nSA, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SDFCHK, nDA_DB_SA, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SDFCHK, nDA_nDB_SA, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SDFCHK, nDA_nDB_nSA, 1'b1);
    tsmc_xbuf (DB_SA_SDFCHK, DB_SA, 1'b1);
    tsmc_xbuf (nDB_SA_SDFCHK, nDB_SA, 1'b1);
    tsmc_xbuf (DA_nSA_SDFCHK, DA_nSA, 1'b1);
    tsmc_xbuf (nDA_nSA_SDFCHK, nDA_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_SDFCHK, DA_nDB, 1'b1);
    tsmc_xbuf (nDA_DB_SDFCHK, nDA_DB, 1'b1);
  `endif

    not (nDA, DA);
    not (nDB, DB);
    not (nSA, SA);
    and (DA_DB_SA, DA, DB, SA);
    and (DA_DB_nSA, DA, DB, nSA);
    and (DA_nDB_SA, DA, nDB, SA);
    and (nDA_DB_nSA, nDA, DB, nSA);
    and (DA_nDB_nSA, DA, nDB, nSA);
    and (nDA_DB_SA, nDA, DB, SA);
    and (nDA_nDB_SA, nDA, nDB, SA);
    and (nDA_nDB_nSA, nDA, nDB, nSA);
    and (DB_SA, DB, SA);
    and (nDB_SA, nDB, SA);
    and (DA_nSA, DA, nSA);
    and (nDA_nSA, nDA, nSA);
    and (DA_nDB, DA, nDB);
    and (nDA_DB, nDA, DB);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SA_int_not, SA_d);
    buf  (DA_check, SA_d);
  `else
    not  (SA_int_not, SA);
    buf  (DA_check, SA);
  `endif
  buf  (DB_check, SA_int_not);
  pullup  (CP_check);
  pullup  (SA_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((DA && DB) || (DA && !(DB) && SA) || (!(DA) && DB && !(SA))))) = (0, 0);
    (posedge CP => (QN-:((DA && DB) || (DA && !(DB) && SA) || (!(DA) && DB && !(SA))))) = (0, 0);
    $width (posedge CP &&& DA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DB_SA_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
  `else
    $setuphold (posedge CP &&& DB_SA_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, negedge SA , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFXQD1 (DA, DB, SA, CP, Q);
    input DA, DB, SA, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire DA_d, DB_d, SA_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB_d, DA_d, SA_d);
        tsmc_dff (Q_buf, D, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB, DA, SA);
        tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (DA_DB_SA_SDFCHK, DA_DB_SA, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SDFCHK, DA_DB_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SDFCHK, DA_nDB_SA, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SDFCHK, nDA_DB_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SDFCHK, DA_nDB_nSA, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SDFCHK, nDA_DB_SA, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SDFCHK, nDA_nDB_SA, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SDFCHK, nDA_nDB_nSA, 1'b1);
    tsmc_xbuf (DB_SA_SDFCHK, DB_SA, 1'b1);
    tsmc_xbuf (nDB_SA_SDFCHK, nDB_SA, 1'b1);
    tsmc_xbuf (DA_nSA_SDFCHK, DA_nSA, 1'b1);
    tsmc_xbuf (nDA_nSA_SDFCHK, nDA_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_SDFCHK, DA_nDB, 1'b1);
    tsmc_xbuf (nDA_DB_SDFCHK, nDA_DB, 1'b1);
  `endif

    not (nDA, DA);
    not (nDB, DB);
    not (nSA, SA);
    and (DA_DB_SA, DA, DB, SA);
    and (DA_DB_nSA, DA, DB, nSA);
    and (DA_nDB_SA, DA, nDB, SA);
    and (nDA_DB_nSA, nDA, DB, nSA);
    and (DA_nDB_nSA, DA, nDB, nSA);
    and (nDA_DB_SA, nDA, DB, SA);
    and (nDA_nDB_SA, nDA, nDB, SA);
    and (nDA_nDB_nSA, nDA, nDB, nSA);
    and (DB_SA, DB, SA);
    and (nDB_SA, nDB, SA);
    and (DA_nSA, DA, nSA);
    and (nDA_nSA, nDA, nSA);
    and (DA_nDB, DA, nDB);
    and (nDA_DB, nDA, DB);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SA_int_not, SA_d);
    buf  (DA_check, SA_d);
  `else
    not  (SA_int_not, SA);
    buf  (DA_check, SA);
  `endif
  buf  (DB_check, SA_int_not);
  pullup  (CP_check);
  pullup  (SA_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((DA && DB) || (DA && !(DB) && SA) || (!(DA) && DB && !(SA))))) = (0, 0);
    $width (posedge CP &&& DA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DB_SA_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
  `else
    $setuphold (posedge CP &&& DB_SA_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, negedge SA , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFXQD2 (DA, DB, SA, CP, Q);
    input DA, DB, SA, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire DA_d, DB_d, SA_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB_d, DA_d, SA_d);
        tsmc_dff (Q_buf, D, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB, DA, SA);
        tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (DA_DB_SA_SDFCHK, DA_DB_SA, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SDFCHK, DA_DB_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SDFCHK, DA_nDB_SA, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SDFCHK, nDA_DB_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SDFCHK, DA_nDB_nSA, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SDFCHK, nDA_DB_SA, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SDFCHK, nDA_nDB_SA, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SDFCHK, nDA_nDB_nSA, 1'b1);
    tsmc_xbuf (DB_SA_SDFCHK, DB_SA, 1'b1);
    tsmc_xbuf (nDB_SA_SDFCHK, nDB_SA, 1'b1);
    tsmc_xbuf (DA_nSA_SDFCHK, DA_nSA, 1'b1);
    tsmc_xbuf (nDA_nSA_SDFCHK, nDA_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_SDFCHK, DA_nDB, 1'b1);
    tsmc_xbuf (nDA_DB_SDFCHK, nDA_DB, 1'b1);
  `endif

    not (nDA, DA);
    not (nDB, DB);
    not (nSA, SA);
    and (DA_DB_SA, DA, DB, SA);
    and (DA_DB_nSA, DA, DB, nSA);
    and (DA_nDB_SA, DA, nDB, SA);
    and (nDA_DB_nSA, nDA, DB, nSA);
    and (DA_nDB_nSA, DA, nDB, nSA);
    and (nDA_DB_SA, nDA, DB, SA);
    and (nDA_nDB_SA, nDA, nDB, SA);
    and (nDA_nDB_nSA, nDA, nDB, nSA);
    and (DB_SA, DB, SA);
    and (nDB_SA, nDB, SA);
    and (DA_nSA, DA, nSA);
    and (nDA_nSA, nDA, nSA);
    and (DA_nDB, DA, nDB);
    and (nDA_DB, nDA, DB);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SA_int_not, SA_d);
    buf  (DA_check, SA_d);
  `else
    not  (SA_int_not, SA);
    buf  (DA_check, SA);
  `endif
  buf  (DB_check, SA_int_not);
  pullup  (CP_check);
  pullup  (SA_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((DA && DB) || (DA && !(DB) && SA) || (!(DA) && DB && !(SA))))) = (0, 0);
    $width (posedge CP &&& DA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DB_SA_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
  `else
    $setuphold (posedge CP &&& DB_SA_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, negedge SA , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFXQD4 (DA, DB, SA, CP, Q);
    input DA, DB, SA, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire DA_d, DB_d, SA_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB_d, DA_d, SA_d);
        tsmc_dff (Q_buf, D, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB, DA, SA);
        tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (DA_DB_SA_SDFCHK, DA_DB_SA, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SDFCHK, DA_DB_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SDFCHK, DA_nDB_SA, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SDFCHK, nDA_DB_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SDFCHK, DA_nDB_nSA, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SDFCHK, nDA_DB_SA, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SDFCHK, nDA_nDB_SA, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SDFCHK, nDA_nDB_nSA, 1'b1);
    tsmc_xbuf (DB_SA_SDFCHK, DB_SA, 1'b1);
    tsmc_xbuf (nDB_SA_SDFCHK, nDB_SA, 1'b1);
    tsmc_xbuf (DA_nSA_SDFCHK, DA_nSA, 1'b1);
    tsmc_xbuf (nDA_nSA_SDFCHK, nDA_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_SDFCHK, DA_nDB, 1'b1);
    tsmc_xbuf (nDA_DB_SDFCHK, nDA_DB, 1'b1);
  `endif

    not (nDA, DA);
    not (nDB, DB);
    not (nSA, SA);
    and (DA_DB_SA, DA, DB, SA);
    and (DA_DB_nSA, DA, DB, nSA);
    and (DA_nDB_SA, DA, nDB, SA);
    and (nDA_DB_nSA, nDA, DB, nSA);
    and (DA_nDB_nSA, DA, nDB, nSA);
    and (nDA_DB_SA, nDA, DB, SA);
    and (nDA_nDB_SA, nDA, nDB, SA);
    and (nDA_nDB_nSA, nDA, nDB, nSA);
    and (DB_SA, DB, SA);
    and (nDB_SA, nDB, SA);
    and (DA_nSA, DA, nSA);
    and (nDA_nSA, nDA, nSA);
    and (DA_nDB, DA, nDB);
    and (nDA_DB, nDA, DB);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SA_int_not, SA_d);
    buf  (DA_check, SA_d);
  `else
    not  (SA_int_not, SA);
    buf  (DA_check, SA);
  `endif
  buf  (DB_check, SA_int_not);
  pullup  (CP_check);
  pullup  (SA_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((DA && DB) || (DA && !(DB) && SA) || (!(DA) && DB && !(SA))))) = (0, 0);
    $width (posedge CP &&& DA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DB_SA_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
  `else
    $setuphold (posedge CP &&& DB_SA_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, negedge SA , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFCND1 (D, E, CP, CDN, Q, QN);
    input D, E, CP, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, E_d, CP_d;
        pullup (SDN);
        tsmc_mux (DE, Q_buf, D_d, E_d);
        tsmc_dff (Q_buf, DE, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (SDN);
        buf (CDN_i, CDN);
        tsmc_mux (DE, Q_buf, D, E);
        tsmc_dff (Q_buf, DE, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_E_SDFCHK, CP_D_E, 1'b1);
    tsmc_xbuf (CP_D_nE_SDFCHK, CP_D_nE, 1'b1);
    tsmc_xbuf (CP_nD_E_SDFCHK, CP_nD_E, 1'b1);
    tsmc_xbuf (CP_nD_nE_SDFCHK, CP_nD_nE, 1'b1);
    tsmc_xbuf (nCP_D_E_SDFCHK, nCP_D_E, 1'b1);
    tsmc_xbuf (nCP_nD_E_SDFCHK, nCP_nD_E, 1'b1);
    tsmc_xbuf (nCP_D_nE_SDFCHK, nCP_D_nE, 1'b1);
    tsmc_xbuf (nCP_nD_nE_SDFCHK, nCP_nD_nE, 1'b1);
    tsmc_xbuf (CDN_D_E_SDFCHK, CDN_D_E, 1'b1);
    tsmc_xbuf (CDN_nD_E_SDFCHK, CDN_nD_E, 1'b1);
    tsmc_xbuf (CDN_E_SDFCHK, CDN_E, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    tsmc_xbuf (D_E_SDFCHK, D_E, 1'b1);
  `endif

    not (nD, D);
    not (nE, E);
    not (nCP, CP);
    and (CP_D_E, CP, D, E);
    and (CP_D_nE, CP, D, nE);
    and (CP_nD_E, CP, nD, E);
    and (CP_nD_nE, CP, nD, nE);
    and (nCP_D_E, nCP, D, E);
    and (nCP_nD_E, nCP, nD, E);
    and (nCP_D_nE, nCP, D, nE);
    and (nCP_nD_nE, nCP, nD, nE);
    and (CDN_D_E, CDN, D, E);
    and (CDN_nD_E, CDN, nD, E);
    and (CDN_E, CDN, E);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);
    and (D_E, D, E);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    and  (D_check, CDN_i, E_d);
  `else
    not  (E_int_not, E);
    and  (D_check, CDN_i, E);
  `endif
  and  (CP_check, CDN_i, D_check);
  buf  (E_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    $width (negedge CDN &&& CP_D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_E_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_D_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $recrem (posedge CDN &&& D_E_SDFCHK, posedge CP &&& D_E_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_E_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_D_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $recovery (posedge CDN &&& D_E_SDFCHK, posedge CP &&& D_E_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_E_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_E_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_E_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDFCHK, negedge E , 0, 0, notifier);
    $recovery (posedge CDN &&& D_E_SDFCHK, posedge CP &&& D_E_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_E_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFCND2 (D, E, CP, CDN, Q, QN);
    input D, E, CP, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, E_d, CP_d;
        pullup (SDN);
        tsmc_mux (DE, Q_buf, D_d, E_d);
        tsmc_dff (Q_buf, DE, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (SDN);
        buf (CDN_i, CDN);
        tsmc_mux (DE, Q_buf, D, E);
        tsmc_dff (Q_buf, DE, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_E_SDFCHK, CP_D_E, 1'b1);
    tsmc_xbuf (CP_D_nE_SDFCHK, CP_D_nE, 1'b1);
    tsmc_xbuf (CP_nD_E_SDFCHK, CP_nD_E, 1'b1);
    tsmc_xbuf (CP_nD_nE_SDFCHK, CP_nD_nE, 1'b1);
    tsmc_xbuf (nCP_D_E_SDFCHK, nCP_D_E, 1'b1);
    tsmc_xbuf (nCP_nD_E_SDFCHK, nCP_nD_E, 1'b1);
    tsmc_xbuf (nCP_D_nE_SDFCHK, nCP_D_nE, 1'b1);
    tsmc_xbuf (nCP_nD_nE_SDFCHK, nCP_nD_nE, 1'b1);
    tsmc_xbuf (CDN_D_E_SDFCHK, CDN_D_E, 1'b1);
    tsmc_xbuf (CDN_nD_E_SDFCHK, CDN_nD_E, 1'b1);
    tsmc_xbuf (CDN_E_SDFCHK, CDN_E, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    tsmc_xbuf (D_E_SDFCHK, D_E, 1'b1);
  `endif

    not (nD, D);
    not (nE, E);
    not (nCP, CP);
    and (CP_D_E, CP, D, E);
    and (CP_D_nE, CP, D, nE);
    and (CP_nD_E, CP, nD, E);
    and (CP_nD_nE, CP, nD, nE);
    and (nCP_D_E, nCP, D, E);
    and (nCP_nD_E, nCP, nD, E);
    and (nCP_D_nE, nCP, D, nE);
    and (nCP_nD_nE, nCP, nD, nE);
    and (CDN_D_E, CDN, D, E);
    and (CDN_nD_E, CDN, nD, E);
    and (CDN_E, CDN, E);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);
    and (D_E, D, E);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    and  (D_check, CDN_i, E_d);
  `else
    not  (E_int_not, E);
    and  (D_check, CDN_i, E);
  `endif
  and  (CP_check, CDN_i, D_check);
  buf  (E_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    $width (negedge CDN &&& CP_D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_E_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_D_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $recrem (posedge CDN &&& D_E_SDFCHK, posedge CP &&& D_E_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_E_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_D_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $recovery (posedge CDN &&& D_E_SDFCHK, posedge CP &&& D_E_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_E_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_E_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_E_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDFCHK, negedge E , 0, 0, notifier);
    $recovery (posedge CDN &&& D_E_SDFCHK, posedge CP &&& D_E_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_E_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFCND4 (D, E, CP, CDN, Q, QN);
    input D, E, CP, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, E_d, CP_d;
        pullup (SDN);
        tsmc_mux (DE, Q_buf, D_d, E_d);
        tsmc_dff (Q_buf, DE, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (SDN);
        buf (CDN_i, CDN);
        tsmc_mux (DE, Q_buf, D, E);
        tsmc_dff (Q_buf, DE, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_E_SDFCHK, CP_D_E, 1'b1);
    tsmc_xbuf (CP_D_nE_SDFCHK, CP_D_nE, 1'b1);
    tsmc_xbuf (CP_nD_E_SDFCHK, CP_nD_E, 1'b1);
    tsmc_xbuf (CP_nD_nE_SDFCHK, CP_nD_nE, 1'b1);
    tsmc_xbuf (nCP_D_E_SDFCHK, nCP_D_E, 1'b1);
    tsmc_xbuf (nCP_nD_E_SDFCHK, nCP_nD_E, 1'b1);
    tsmc_xbuf (nCP_D_nE_SDFCHK, nCP_D_nE, 1'b1);
    tsmc_xbuf (nCP_nD_nE_SDFCHK, nCP_nD_nE, 1'b1);
    tsmc_xbuf (CDN_D_E_SDFCHK, CDN_D_E, 1'b1);
    tsmc_xbuf (CDN_nD_E_SDFCHK, CDN_nD_E, 1'b1);
    tsmc_xbuf (CDN_E_SDFCHK, CDN_E, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    tsmc_xbuf (D_E_SDFCHK, D_E, 1'b1);
  `endif

    not (nD, D);
    not (nE, E);
    not (nCP, CP);
    and (CP_D_E, CP, D, E);
    and (CP_D_nE, CP, D, nE);
    and (CP_nD_E, CP, nD, E);
    and (CP_nD_nE, CP, nD, nE);
    and (nCP_D_E, nCP, D, E);
    and (nCP_nD_E, nCP, nD, E);
    and (nCP_D_nE, nCP, D, nE);
    and (nCP_nD_nE, nCP, nD, nE);
    and (CDN_D_E, CDN, D, E);
    and (CDN_nD_E, CDN, nD, E);
    and (CDN_E, CDN, E);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);
    and (D_E, D, E);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    and  (D_check, CDN_i, E_d);
  `else
    not  (E_int_not, E);
    and  (D_check, CDN_i, E);
  `endif
  and  (CP_check, CDN_i, D_check);
  buf  (E_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    $width (negedge CDN &&& CP_D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_E_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_D_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $recrem (posedge CDN &&& D_E_SDFCHK, posedge CP &&& D_E_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_E_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_D_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $recovery (posedge CDN &&& D_E_SDFCHK, posedge CP &&& D_E_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_E_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_E_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_E_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDFCHK, negedge E , 0, 0, notifier);
    $recovery (posedge CDN &&& D_E_SDFCHK, posedge CP &&& D_E_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_E_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFCNQD1 (D, E, CP, CDN, Q);
    input D, E, CP, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, E_d, CP_d;
        pullup (SDN);
        tsmc_mux (DE, Q_buf, D_d, E_d);
        tsmc_dff (Q_buf, DE, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (SDN);
        buf (CDN_i, CDN);
        tsmc_mux (DE, Q_buf, D, E);
        tsmc_dff (Q_buf, DE, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_E_SDFCHK, CP_D_E, 1'b1);
    tsmc_xbuf (CP_D_nE_SDFCHK, CP_D_nE, 1'b1);
    tsmc_xbuf (CP_nD_E_SDFCHK, CP_nD_E, 1'b1);
    tsmc_xbuf (CP_nD_nE_SDFCHK, CP_nD_nE, 1'b1);
    tsmc_xbuf (nCP_D_E_SDFCHK, nCP_D_E, 1'b1);
    tsmc_xbuf (nCP_nD_E_SDFCHK, nCP_nD_E, 1'b1);
    tsmc_xbuf (nCP_D_nE_SDFCHK, nCP_D_nE, 1'b1);
    tsmc_xbuf (nCP_nD_nE_SDFCHK, nCP_nD_nE, 1'b1);
    tsmc_xbuf (CDN_D_E_SDFCHK, CDN_D_E, 1'b1);
    tsmc_xbuf (CDN_nD_E_SDFCHK, CDN_nD_E, 1'b1);
    tsmc_xbuf (CDN_E_SDFCHK, CDN_E, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    tsmc_xbuf (D_E_SDFCHK, D_E, 1'b1);
  `endif

    not (nD, D);
    not (nE, E);
    not (nCP, CP);
    and (CP_D_E, CP, D, E);
    and (CP_D_nE, CP, D, nE);
    and (CP_nD_E, CP, nD, E);
    and (CP_nD_nE, CP, nD, nE);
    and (nCP_D_E, nCP, D, E);
    and (nCP_nD_E, nCP, nD, E);
    and (nCP_D_nE, nCP, D, nE);
    and (nCP_nD_nE, nCP, nD, nE);
    and (CDN_D_E, CDN, D, E);
    and (CDN_nD_E, CDN, nD, E);
    and (CDN_E, CDN, E);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);
    and (D_E, D, E);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    and  (D_check, CDN_i, E_d);
  `else
    not  (E_int_not, E);
    and  (D_check, CDN_i, E);
  `endif
  and  (CP_check, CDN_i, D_check);
  buf  (E_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    $width (negedge CDN &&& CP_D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_E_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_D_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $recrem (posedge CDN &&& D_E_SDFCHK, posedge CP &&& D_E_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_E_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_D_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $recovery (posedge CDN &&& D_E_SDFCHK, posedge CP &&& D_E_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_E_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_E_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_E_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDFCHK, negedge E , 0, 0, notifier);
    $recovery (posedge CDN &&& D_E_SDFCHK, posedge CP &&& D_E_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_E_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFCNQD2 (D, E, CP, CDN, Q);
    input D, E, CP, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, E_d, CP_d;
        pullup (SDN);
        tsmc_mux (DE, Q_buf, D_d, E_d);
        tsmc_dff (Q_buf, DE, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (SDN);
        buf (CDN_i, CDN);
        tsmc_mux (DE, Q_buf, D, E);
        tsmc_dff (Q_buf, DE, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_E_SDFCHK, CP_D_E, 1'b1);
    tsmc_xbuf (CP_D_nE_SDFCHK, CP_D_nE, 1'b1);
    tsmc_xbuf (CP_nD_E_SDFCHK, CP_nD_E, 1'b1);
    tsmc_xbuf (CP_nD_nE_SDFCHK, CP_nD_nE, 1'b1);
    tsmc_xbuf (nCP_D_E_SDFCHK, nCP_D_E, 1'b1);
    tsmc_xbuf (nCP_nD_E_SDFCHK, nCP_nD_E, 1'b1);
    tsmc_xbuf (nCP_D_nE_SDFCHK, nCP_D_nE, 1'b1);
    tsmc_xbuf (nCP_nD_nE_SDFCHK, nCP_nD_nE, 1'b1);
    tsmc_xbuf (CDN_D_E_SDFCHK, CDN_D_E, 1'b1);
    tsmc_xbuf (CDN_nD_E_SDFCHK, CDN_nD_E, 1'b1);
    tsmc_xbuf (CDN_E_SDFCHK, CDN_E, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    tsmc_xbuf (D_E_SDFCHK, D_E, 1'b1);
  `endif

    not (nD, D);
    not (nE, E);
    not (nCP, CP);
    and (CP_D_E, CP, D, E);
    and (CP_D_nE, CP, D, nE);
    and (CP_nD_E, CP, nD, E);
    and (CP_nD_nE, CP, nD, nE);
    and (nCP_D_E, nCP, D, E);
    and (nCP_nD_E, nCP, nD, E);
    and (nCP_D_nE, nCP, D, nE);
    and (nCP_nD_nE, nCP, nD, nE);
    and (CDN_D_E, CDN, D, E);
    and (CDN_nD_E, CDN, nD, E);
    and (CDN_E, CDN, E);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);
    and (D_E, D, E);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    and  (D_check, CDN_i, E_d);
  `else
    not  (E_int_not, E);
    and  (D_check, CDN_i, E);
  `endif
  and  (CP_check, CDN_i, D_check);
  buf  (E_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    $width (negedge CDN &&& CP_D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_E_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_D_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $recrem (posedge CDN &&& D_E_SDFCHK, posedge CP &&& D_E_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_E_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_D_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $recovery (posedge CDN &&& D_E_SDFCHK, posedge CP &&& D_E_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_E_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_E_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_E_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDFCHK, negedge E , 0, 0, notifier);
    $recovery (posedge CDN &&& D_E_SDFCHK, posedge CP &&& D_E_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_E_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFCNQD4 (D, E, CP, CDN, Q);
    input D, E, CP, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, E_d, CP_d;
        pullup (SDN);
        tsmc_mux (DE, Q_buf, D_d, E_d);
        tsmc_dff (Q_buf, DE, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (SDN);
        buf (CDN_i, CDN);
        tsmc_mux (DE, Q_buf, D, E);
        tsmc_dff (Q_buf, DE, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_E_SDFCHK, CP_D_E, 1'b1);
    tsmc_xbuf (CP_D_nE_SDFCHK, CP_D_nE, 1'b1);
    tsmc_xbuf (CP_nD_E_SDFCHK, CP_nD_E, 1'b1);
    tsmc_xbuf (CP_nD_nE_SDFCHK, CP_nD_nE, 1'b1);
    tsmc_xbuf (nCP_D_E_SDFCHK, nCP_D_E, 1'b1);
    tsmc_xbuf (nCP_nD_E_SDFCHK, nCP_nD_E, 1'b1);
    tsmc_xbuf (nCP_D_nE_SDFCHK, nCP_D_nE, 1'b1);
    tsmc_xbuf (nCP_nD_nE_SDFCHK, nCP_nD_nE, 1'b1);
    tsmc_xbuf (CDN_D_E_SDFCHK, CDN_D_E, 1'b1);
    tsmc_xbuf (CDN_nD_E_SDFCHK, CDN_nD_E, 1'b1);
    tsmc_xbuf (CDN_E_SDFCHK, CDN_E, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    tsmc_xbuf (D_E_SDFCHK, D_E, 1'b1);
  `endif

    not (nD, D);
    not (nE, E);
    not (nCP, CP);
    and (CP_D_E, CP, D, E);
    and (CP_D_nE, CP, D, nE);
    and (CP_nD_E, CP, nD, E);
    and (CP_nD_nE, CP, nD, nE);
    and (nCP_D_E, nCP, D, E);
    and (nCP_nD_E, nCP, nD, E);
    and (nCP_D_nE, nCP, D, nE);
    and (nCP_nD_nE, nCP, nD, nE);
    and (CDN_D_E, CDN, D, E);
    and (CDN_nD_E, CDN, nD, E);
    and (CDN_E, CDN, E);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);
    and (D_E, D, E);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    and  (D_check, CDN_i, E_d);
  `else
    not  (E_int_not, E);
    and  (D_check, CDN_i, E);
  `endif
  and  (CP_check, CDN_i, D_check);
  buf  (E_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    $width (negedge CDN &&& CP_D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_E_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_D_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $recrem (posedge CDN &&& D_E_SDFCHK, posedge CP &&& D_E_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_E_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_D_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $recovery (posedge CDN &&& D_E_SDFCHK, posedge CP &&& D_E_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_E_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_E_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_E_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDFCHK, negedge E , 0, 0, notifier);
    $recovery (posedge CDN &&& D_E_SDFCHK, posedge CP &&& D_E_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_E_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFD1 (D, E, CP, Q, QN);
    input D, E, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, E_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (DE, Q_buf, D_d, E_d);
        tsmc_dff (Q_buf, DE, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (DE, Q_buf, D, E);
        tsmc_dff (Q_buf, DE, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_SDFCHK, E, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_E_SDFCHK, D_E, 1'b1);
    tsmc_xbuf (nD_E_SDFCHK, nD_E, 1'b1);
  `endif

    not (nD, D);
    and (D_E, D, E);
    and (nD_E, nD, E);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    buf  (D_check, E_d);
  `else
    not  (E_int_not, E);
    buf  (D_check, E);
  `endif
  buf  (CP_check, D_check);
  pullup  (E_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    (posedge CP => (QN-:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& E_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
  `else
    $setuphold (posedge CP &&& E_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDFCHK, negedge E , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFD2 (D, E, CP, Q, QN);
    input D, E, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, E_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (DE, Q_buf, D_d, E_d);
        tsmc_dff (Q_buf, DE, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (DE, Q_buf, D, E);
        tsmc_dff (Q_buf, DE, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_SDFCHK, E, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_E_SDFCHK, D_E, 1'b1);
    tsmc_xbuf (nD_E_SDFCHK, nD_E, 1'b1);
  `endif

    not (nD, D);
    and (D_E, D, E);
    and (nD_E, nD, E);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    buf  (D_check, E_d);
  `else
    not  (E_int_not, E);
    buf  (D_check, E);
  `endif
  buf  (CP_check, D_check);
  pullup  (E_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    (posedge CP => (QN-:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& E_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
  `else
    $setuphold (posedge CP &&& E_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDFCHK, negedge E , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFD4 (D, E, CP, Q, QN);
    input D, E, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, E_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (DE, Q_buf, D_d, E_d);
        tsmc_dff (Q_buf, DE, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (DE, Q_buf, D, E);
        tsmc_dff (Q_buf, DE, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_SDFCHK, E, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_E_SDFCHK, D_E, 1'b1);
    tsmc_xbuf (nD_E_SDFCHK, nD_E, 1'b1);
  `endif

    not (nD, D);
    and (D_E, D, E);
    and (nD_E, nD, E);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    buf  (D_check, E_d);
  `else
    not  (E_int_not, E);
    buf  (D_check, E);
  `endif
  buf  (CP_check, D_check);
  pullup  (E_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    (posedge CP => (QN-:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& E_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
  `else
    $setuphold (posedge CP &&& E_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDFCHK, negedge E , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFKCND1 (D, E, CP, CN, Q, QN);
    input D, E, CP, CN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, E_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        and (D2, CN_d, D1);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        and (D2, CN, D1);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_E_SDFCHK, CN_D_E, 1'b1);
    tsmc_xbuf (CN_nD_E_SDFCHK, CN_nD_E, 1'b1);
    tsmc_xbuf (nCN_D_E_SDFCHK, nCN_D_E, 1'b1);
    tsmc_xbuf (nCN_D_nE_SDFCHK, nCN_D_nE, 1'b1);
    tsmc_xbuf (nCN_nD_E_SDFCHK, nCN_nD_E, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SDFCHK, nCN_nD_nE, 1'b1);
    tsmc_xbuf (D_E_SDFCHK, D_E, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    tsmc_xbuf (CN_E_SDFCHK, CN_E, 1'b1);
    tsmc_xbuf (CN_D_SDFCHK, CN_D, 1'b1);
    tsmc_xbuf (CN_nD_SDFCHK, CN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nE, E);
    not (nCN, CN);
    and (CN_D_E, CN, D, E);
    and (CN_nD_E, CN, nD, E);
    and (nCN_D_E, nCN, D, E);
    and (nCN_D_nE, nCN, D, nE);
    and (nCN_nD_E, nCN, nD, E);
    and (nCN_nD_nE, nCN, nD, nE);
    and (D_E, D, E);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);
    and (CN_E, CN, E);
    and (CN_D, CN, D);
    and (CN_nD, CN, nD);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (CN_int_not, CN_d);
    buf  (E_check, CN_d);
    and  (D_check, CN_d, E_d);
  `else
    not  (CN_int_not, CN);
    buf  (E_check, CN);
    and  (D_check, CN, E);
  `endif
  or   (CP_check, CN_int_not, D_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((CN && E && D) || (CN && !(E) && Q_buf)))) = (0, 0);
    (posedge CP => (QN-:((CN && E && D) || (CN && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CN_D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_E_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_E_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_E_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_E_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_D_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
  `else
    $setuphold (posedge CP &&& D_E_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, negedge E , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFKCND2 (D, E, CP, CN, Q, QN);
    input D, E, CP, CN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, E_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        and (D2, CN_d, D1);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        and (D2, CN, D1);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_E_SDFCHK, CN_D_E, 1'b1);
    tsmc_xbuf (CN_nD_E_SDFCHK, CN_nD_E, 1'b1);
    tsmc_xbuf (nCN_D_E_SDFCHK, nCN_D_E, 1'b1);
    tsmc_xbuf (nCN_D_nE_SDFCHK, nCN_D_nE, 1'b1);
    tsmc_xbuf (nCN_nD_E_SDFCHK, nCN_nD_E, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SDFCHK, nCN_nD_nE, 1'b1);
    tsmc_xbuf (D_E_SDFCHK, D_E, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    tsmc_xbuf (CN_E_SDFCHK, CN_E, 1'b1);
    tsmc_xbuf (CN_D_SDFCHK, CN_D, 1'b1);
    tsmc_xbuf (CN_nD_SDFCHK, CN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nE, E);
    not (nCN, CN);
    and (CN_D_E, CN, D, E);
    and (CN_nD_E, CN, nD, E);
    and (nCN_D_E, nCN, D, E);
    and (nCN_D_nE, nCN, D, nE);
    and (nCN_nD_E, nCN, nD, E);
    and (nCN_nD_nE, nCN, nD, nE);
    and (D_E, D, E);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);
    and (CN_E, CN, E);
    and (CN_D, CN, D);
    and (CN_nD, CN, nD);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (CN_int_not, CN_d);
    buf  (E_check, CN_d);
    and  (D_check, CN_d, E_d);
  `else
    not  (CN_int_not, CN);
    buf  (E_check, CN);
    and  (D_check, CN, E);
  `endif
  or   (CP_check, CN_int_not, D_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((CN && E && D) || (CN && !(E) && Q_buf)))) = (0, 0);
    (posedge CP => (QN-:((CN && E && D) || (CN && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CN_D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_E_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_E_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_E_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_E_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_D_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
  `else
    $setuphold (posedge CP &&& D_E_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, negedge E , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFKCND4 (D, E, CP, CN, Q, QN);
    input D, E, CP, CN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, E_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        and (D2, CN_d, D1);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        and (D2, CN, D1);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_E_SDFCHK, CN_D_E, 1'b1);
    tsmc_xbuf (CN_nD_E_SDFCHK, CN_nD_E, 1'b1);
    tsmc_xbuf (nCN_D_E_SDFCHK, nCN_D_E, 1'b1);
    tsmc_xbuf (nCN_D_nE_SDFCHK, nCN_D_nE, 1'b1);
    tsmc_xbuf (nCN_nD_E_SDFCHK, nCN_nD_E, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SDFCHK, nCN_nD_nE, 1'b1);
    tsmc_xbuf (D_E_SDFCHK, D_E, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    tsmc_xbuf (CN_E_SDFCHK, CN_E, 1'b1);
    tsmc_xbuf (CN_D_SDFCHK, CN_D, 1'b1);
    tsmc_xbuf (CN_nD_SDFCHK, CN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nE, E);
    not (nCN, CN);
    and (CN_D_E, CN, D, E);
    and (CN_nD_E, CN, nD, E);
    and (nCN_D_E, nCN, D, E);
    and (nCN_D_nE, nCN, D, nE);
    and (nCN_nD_E, nCN, nD, E);
    and (nCN_nD_nE, nCN, nD, nE);
    and (D_E, D, E);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);
    and (CN_E, CN, E);
    and (CN_D, CN, D);
    and (CN_nD, CN, nD);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (CN_int_not, CN_d);
    buf  (E_check, CN_d);
    and  (D_check, CN_d, E_d);
  `else
    not  (CN_int_not, CN);
    buf  (E_check, CN);
    and  (D_check, CN, E);
  `endif
  or   (CP_check, CN_int_not, D_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((CN && E && D) || (CN && !(E) && Q_buf)))) = (0, 0);
    (posedge CP => (QN-:((CN && E && D) || (CN && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CN_D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_E_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_E_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_E_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_E_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_D_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
  `else
    $setuphold (posedge CP &&& D_E_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, negedge E , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFKCNQD1 (D, E, CP, CN, Q);
    input D, E, CP, CN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire D_d, E_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        and (D2, CN_d, D1);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        and (D2, CN, D1);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_E_SDFCHK, CN_D_E, 1'b1);
    tsmc_xbuf (CN_nD_E_SDFCHK, CN_nD_E, 1'b1);
    tsmc_xbuf (nCN_D_E_SDFCHK, nCN_D_E, 1'b1);
    tsmc_xbuf (nCN_D_nE_SDFCHK, nCN_D_nE, 1'b1);
    tsmc_xbuf (nCN_nD_E_SDFCHK, nCN_nD_E, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SDFCHK, nCN_nD_nE, 1'b1);
    tsmc_xbuf (D_E_SDFCHK, D_E, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    tsmc_xbuf (CN_E_SDFCHK, CN_E, 1'b1);
    tsmc_xbuf (CN_D_SDFCHK, CN_D, 1'b1);
    tsmc_xbuf (CN_nD_SDFCHK, CN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nE, E);
    not (nCN, CN);
    and (CN_D_E, CN, D, E);
    and (CN_nD_E, CN, nD, E);
    and (nCN_D_E, nCN, D, E);
    and (nCN_D_nE, nCN, D, nE);
    and (nCN_nD_E, nCN, nD, E);
    and (nCN_nD_nE, nCN, nD, nE);
    and (D_E, D, E);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);
    and (CN_E, CN, E);
    and (CN_D, CN, D);
    and (CN_nD, CN, nD);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (CN_int_not, CN_d);
    buf  (E_check, CN_d);
    and  (D_check, CN_d, E_d);
  `else
    not  (CN_int_not, CN);
    buf  (E_check, CN);
    and  (D_check, CN, E);
  `endif
  or   (CP_check, CN_int_not, D_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((CN && E && D) || (CN && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CN_D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_E_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_E_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_E_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_E_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_D_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
  `else
    $setuphold (posedge CP &&& D_E_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, negedge E , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFKCNQD2 (D, E, CP, CN, Q);
    input D, E, CP, CN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire D_d, E_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        and (D2, CN_d, D1);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        and (D2, CN, D1);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_E_SDFCHK, CN_D_E, 1'b1);
    tsmc_xbuf (CN_nD_E_SDFCHK, CN_nD_E, 1'b1);
    tsmc_xbuf (nCN_D_E_SDFCHK, nCN_D_E, 1'b1);
    tsmc_xbuf (nCN_D_nE_SDFCHK, nCN_D_nE, 1'b1);
    tsmc_xbuf (nCN_nD_E_SDFCHK, nCN_nD_E, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SDFCHK, nCN_nD_nE, 1'b1);
    tsmc_xbuf (D_E_SDFCHK, D_E, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    tsmc_xbuf (CN_E_SDFCHK, CN_E, 1'b1);
    tsmc_xbuf (CN_D_SDFCHK, CN_D, 1'b1);
    tsmc_xbuf (CN_nD_SDFCHK, CN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nE, E);
    not (nCN, CN);
    and (CN_D_E, CN, D, E);
    and (CN_nD_E, CN, nD, E);
    and (nCN_D_E, nCN, D, E);
    and (nCN_D_nE, nCN, D, nE);
    and (nCN_nD_E, nCN, nD, E);
    and (nCN_nD_nE, nCN, nD, nE);
    and (D_E, D, E);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);
    and (CN_E, CN, E);
    and (CN_D, CN, D);
    and (CN_nD, CN, nD);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (CN_int_not, CN_d);
    buf  (E_check, CN_d);
    and  (D_check, CN_d, E_d);
  `else
    not  (CN_int_not, CN);
    buf  (E_check, CN);
    and  (D_check, CN, E);
  `endif
  or   (CP_check, CN_int_not, D_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((CN && E && D) || (CN && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CN_D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_E_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_E_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_E_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_E_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_D_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
  `else
    $setuphold (posedge CP &&& D_E_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, negedge E , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFKCNQD4 (D, E, CP, CN, Q);
    input D, E, CP, CN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire D_d, E_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        and (D2, CN_d, D1);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        and (D2, CN, D1);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_E_SDFCHK, CN_D_E, 1'b1);
    tsmc_xbuf (CN_nD_E_SDFCHK, CN_nD_E, 1'b1);
    tsmc_xbuf (nCN_D_E_SDFCHK, nCN_D_E, 1'b1);
    tsmc_xbuf (nCN_D_nE_SDFCHK, nCN_D_nE, 1'b1);
    tsmc_xbuf (nCN_nD_E_SDFCHK, nCN_nD_E, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SDFCHK, nCN_nD_nE, 1'b1);
    tsmc_xbuf (D_E_SDFCHK, D_E, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    tsmc_xbuf (CN_E_SDFCHK, CN_E, 1'b1);
    tsmc_xbuf (CN_D_SDFCHK, CN_D, 1'b1);
    tsmc_xbuf (CN_nD_SDFCHK, CN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nE, E);
    not (nCN, CN);
    and (CN_D_E, CN, D, E);
    and (CN_nD_E, CN, nD, E);
    and (nCN_D_E, nCN, D, E);
    and (nCN_D_nE, nCN, D, nE);
    and (nCN_nD_E, nCN, nD, E);
    and (nCN_nD_nE, nCN, nD, nE);
    and (D_E, D, E);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);
    and (CN_E, CN, E);
    and (CN_D, CN, D);
    and (CN_nD, CN, nD);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (CN_int_not, CN_d);
    buf  (E_check, CN_d);
    and  (D_check, CN_d, E_d);
  `else
    not  (CN_int_not, CN);
    buf  (E_check, CN);
    and  (D_check, CN, E);
  `endif
  or   (CP_check, CN_int_not, D_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((CN && E && D) || (CN && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CN_D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_E_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_E_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_E_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_E_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_D_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
  `else
    $setuphold (posedge CP &&& D_E_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, negedge E , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFQD1 (D, E, CP, Q);
    input D, E, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire D_d, E_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (DE, Q_buf, D_d, E_d);
        tsmc_dff (Q_buf, DE, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (DE, Q_buf, D, E);
        tsmc_dff (Q_buf, DE, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_SDFCHK, E, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_E_SDFCHK, D_E, 1'b1);
    tsmc_xbuf (nD_E_SDFCHK, nD_E, 1'b1);
  `endif

    not (nD, D);
    and (D_E, D, E);
    and (nD_E, nD, E);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    buf  (D_check, E_d);
  `else
    not  (E_int_not, E);
    buf  (D_check, E);
  `endif
  buf  (CP_check, D_check);
  pullup  (E_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& E_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
  `else
    $setuphold (posedge CP &&& E_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDFCHK, negedge E , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFQD2 (D, E, CP, Q);
    input D, E, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire D_d, E_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (DE, Q_buf, D_d, E_d);
        tsmc_dff (Q_buf, DE, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (DE, Q_buf, D, E);
        tsmc_dff (Q_buf, DE, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_SDFCHK, E, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_E_SDFCHK, D_E, 1'b1);
    tsmc_xbuf (nD_E_SDFCHK, nD_E, 1'b1);
  `endif

    not (nD, D);
    and (D_E, D, E);
    and (nD_E, nD, E);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    buf  (D_check, E_d);
  `else
    not  (E_int_not, E);
    buf  (D_check, E);
  `endif
  buf  (CP_check, D_check);
  pullup  (E_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& E_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
  `else
    $setuphold (posedge CP &&& E_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDFCHK, negedge E , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFQD4 (D, E, CP, Q);
    input D, E, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire D_d, E_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (DE, Q_buf, D_d, E_d);
        tsmc_dff (Q_buf, DE, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (DE, Q_buf, D, E);
        tsmc_dff (Q_buf, DE, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_SDFCHK, E, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_E_SDFCHK, D_E, 1'b1);
    tsmc_xbuf (nD_E_SDFCHK, nD_E, 1'b1);
  `endif

    not (nD, D);
    and (D_E, D, E);
    and (nD_E, nD, E);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    buf  (D_check, E_d);
  `else
    not  (E_int_not, E);
    buf  (D_check, E);
  `endif
  buf  (CP_check, D_check);
  pullup  (E_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& D_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& E_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
  `else
    $setuphold (posedge CP &&& E_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDFCHK, negedge E , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module FA1D0 (A, B, CI, S, CO);
    input A, B, CI;
    output S, CO;
    xor (I0_out, A, B);
    xor (S, I0_out, CI);
    and (I1_out, A, B);
    and (I2_out, B, CI);
    and (I3_out, A, CI);
    or (CO, I1_out, I2_out, I3_out);

  specify
    if (B == 1'b1 && CI == 1'b0)
    (A => CO) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => CO) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => CO) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => CO) = (0, 0);
    if (B == 1'b1 && CI == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1)
    (CI => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FA1D1 (A, B, CI, S, CO);
    input A, B, CI;
    output S, CO;
    xor (I0_out, A, B);
    xor (S, I0_out, CI);
    and (I1_out, A, B);
    and (I2_out, B, CI);
    and (I3_out, A, CI);
    or (CO, I1_out, I2_out, I3_out);

  specify
    if (B == 1'b1 && CI == 1'b0)
    (A => CO) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => CO) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => CO) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => CO) = (0, 0);
    if (B == 1'b1 && CI == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1)
    (CI => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FA1D2 (A, B, CI, S, CO);
    input A, B, CI;
    output S, CO;
    xor (I0_out, A, B);
    xor (S, I0_out, CI);
    and (I1_out, A, B);
    and (I2_out, B, CI);
    and (I3_out, A, CI);
    or (CO, I1_out, I2_out, I3_out);

  specify
    if (B == 1'b1 && CI == 1'b0)
    (A => CO) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => CO) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => CO) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => CO) = (0, 0);
    if (B == 1'b1 && CI == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1)
    (CI => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FA1D4 (A, B, CI, S, CO);
    input A, B, CI;
    output S, CO;
    xor (I0_out, A, B);
    xor (S, I0_out, CI);
    and (I1_out, A, B);
    and (I2_out, B, CI);
    and (I3_out, A, CI);
    or (CO, I1_out, I2_out, I3_out);

  specify
    if (B == 1'b1 && CI == 1'b0)
    (A => CO) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => CO) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => CO) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => CO) = (0, 0);
    if (B == 1'b1 && CI == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1)
    (CI => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FCICIND1 (A, B, CIN, CO);
    input A, B, CIN;
    output CO;
    not (I0_out, CIN);
    and (I1_out, I0_out, A);
    and (I2_out, A, B);
    not (I3_out, CIN);
    and (I4_out, B, I3_out);
    or (CO, I1_out, I2_out, I4_out);

  specify
    if (B == 1'b1 && CIN == 1'b1)
    (A => CO) = (0, 0);
    if (B == 1'b0 && CIN == 1'b0)
    (A => CO) = (0, 0);
    if (A == 1'b1 && CIN == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b0 && CIN == 1'b0)
    (B => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CIN => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CIN => CO) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FCICIND2 (A, B, CIN, CO);
    input A, B, CIN;
    output CO;
    not (I0_out, CIN);
    and (I1_out, I0_out, A);
    and (I2_out, A, B);
    not (I3_out, CIN);
    and (I4_out, B, I3_out);
    or (CO, I1_out, I2_out, I4_out);

  specify
    if (B == 1'b1 && CIN == 1'b1)
    (A => CO) = (0, 0);
    if (B == 1'b0 && CIN == 1'b0)
    (A => CO) = (0, 0);
    if (A == 1'b1 && CIN == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b0 && CIN == 1'b0)
    (B => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CIN => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CIN => CO) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FCICOND1 (A, B, CI, CON);
    input A, B, CI;
    output CON;
    and (I0_out, A, B);
    and (I1_out, B, CI);
    and (I2_out, CI, A);
    or (I3_out, I0_out, I1_out, I2_out);
    not (CON, I3_out);

  specify
    if (B == 1'b1 && CI == 1'b0)
    (A => CON) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => CON) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => CON) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => CON) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => CON) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => CON) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FCICOND2 (A, B, CI, CON);
    input A, B, CI;
    output CON;
    and (I0_out, A, B);
    and (I1_out, B, CI);
    and (I2_out, CI, A);
    or (I3_out, I0_out, I1_out, I2_out);
    not (CON, I3_out);

  specify
    if (B == 1'b1 && CI == 1'b0)
    (A => CON) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => CON) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => CON) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => CON) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => CON) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => CON) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FCSICIND1 (A, B, CIN0, CIN1, CS, S, CO0, CO1);
    input A, B, CIN0, CIN1, CS;
    output S, CO0, CO1;
    tsmc_mux (I0_out, CIN0, CIN1, CS);
    xor (I1_out, I0_out, A);
    xor (I2_out, I1_out, B);
    not (S, I2_out);
    not (I4_out, B);
    not (I5_out, A);
    and (I6_out, I4_out, I5_out);
    not (I7_out, A);
    and (I8_out, I7_out, CIN0);
    not (I10_out, B);
    and (I11_out, CIN0, I10_out);
    or (I12_out, I6_out, I8_out, I11_out);
    not (CO0, I12_out);
    not (I14_out, B);
    not (I15_out, A);
    and (I16_out, I14_out, I15_out);
    not (I17_out, A);
    and (I18_out, I17_out, CIN1);
    not (I20_out, B);
    and (I21_out, CIN1, I20_out);
    or (I22_out, I16_out, I18_out, I21_out);
    not (CO1, I22_out);

  specify
    if (B == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b1)
    (A => CO0) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b0)
    (A => CO0) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b1)
    (A => CO0) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b0)
    (A => CO0) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b1)
    (A => CO0) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b0)
    (A => CO0) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b1)
    (A => CO0) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b0)
    (A => CO0) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b1)
    (B => CO0) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b0)
    (B => CO0) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b1)
    (B => CO0) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b0)
    (B => CO0) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b1)
    (B => CO0) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b0)
    (B => CO0) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b1)
    (B => CO0) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b0)
    (B => CO0) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN1 == 1'b1 && CS == 1'b1)
    (CIN0 => CO0) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN1 == 1'b0 && CS == 1'b1)
    (CIN0 => CO0) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN1 == 1'b1 && CS == 1'b1)
    (CIN0 => CO0) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN1 == 1'b0 && CS == 1'b1)
    (CIN0 => CO0) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN1 == 1'b1 && CS == 1'b0)
    (CIN0 => CO0) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN1 == 1'b0 && CS == 1'b0)
    (CIN0 => CO0) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN1 == 1'b1 && CS == 1'b0)
    (CIN0 => CO0) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN1 == 1'b0 && CS == 1'b0)
    (CIN0 => CO0) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b1)
    (A => CO1) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b0)
    (A => CO1) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b1)
    (A => CO1) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b0)
    (A => CO1) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b1)
    (A => CO1) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b0)
    (A => CO1) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b1)
    (A => CO1) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b0)
    (A => CO1) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b1)
    (B => CO1) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b0)
    (B => CO1) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b1)
    (B => CO1) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b0)
    (B => CO1) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b1)
    (B => CO1) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b0)
    (B => CO1) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b1)
    (B => CO1) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b0)
    (B => CO1) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN0 == 1'b1 && CS == 1'b1)
    (CIN1 => CO1) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN0 == 1'b0 && CS == 1'b1)
    (CIN1 => CO1) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN0 == 1'b1 && CS == 1'b1)
    (CIN1 => CO1) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN0 == 1'b0 && CS == 1'b1)
    (CIN1 => CO1) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN0 == 1'b1 && CS == 1'b0)
    (CIN1 => CO1) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN0 == 1'b0 && CS == 1'b0)
    (CIN1 => CO1) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN0 == 1'b1 && CS == 1'b0)
    (CIN1 => CO1) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN0 == 1'b0 && CS == 1'b0)
    (CIN1 => CO1) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN1 == 1'b1 && CS == 1'b0)
    (CIN0 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN1 == 1'b0 && CS == 1'b0)
    (CIN0 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN1 == 1'b1 && CS == 1'b0)
    (CIN0 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN1 == 1'b0 && CS == 1'b0)
    (CIN0 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIN1 == 1'b1 && CS == 1'b0)
    (CIN0 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIN1 == 1'b0 && CS == 1'b0)
    (CIN0 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIN1 == 1'b1 && CS == 1'b0)
    (CIN0 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIN1 == 1'b0 && CS == 1'b0)
    (CIN0 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN0 == 1'b1 && CS == 1'b1)
    (CIN1 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN0 == 1'b0 && CS == 1'b1)
    (CIN1 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN0 == 1'b1 && CS == 1'b1)
    (CIN1 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN0 == 1'b0 && CS == 1'b1)
    (CIN1 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIN0 == 1'b1 && CS == 1'b1)
    (CIN1 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIN0 == 1'b0 && CS == 1'b1)
    (CIN1 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIN0 == 1'b1 && CS == 1'b1)
    (CIN1 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIN0 == 1'b0 && CS == 1'b1)
    (CIN1 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b0)
    (CS => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b0)
    (CS => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b1)
    (CS => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b1)
    (CS => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b1)
    (CS => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b1)
    (CS => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b0)
    (CS => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b0)
    (CS => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FCSICIND2 (A, B, CIN0, CIN1, CS, S, CO0, CO1);
    input A, B, CIN0, CIN1, CS;
    output S, CO0, CO1;
    tsmc_mux (I0_out, CIN0, CIN1, CS);
    xor (I1_out, I0_out, A);
    xor (I2_out, I1_out, B);
    not (S, I2_out);
    not (I4_out, B);
    not (I5_out, A);
    and (I6_out, I4_out, I5_out);
    not (I7_out, A);
    and (I8_out, I7_out, CIN0);
    not (I10_out, B);
    and (I11_out, CIN0, I10_out);
    or (I12_out, I6_out, I8_out, I11_out);
    not (CO0, I12_out);
    not (I14_out, B);
    not (I15_out, A);
    and (I16_out, I14_out, I15_out);
    not (I17_out, A);
    and (I18_out, I17_out, CIN1);
    not (I20_out, B);
    and (I21_out, CIN1, I20_out);
    or (I22_out, I16_out, I18_out, I21_out);
    not (CO1, I22_out);

  specify
    if (B == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b1)
    (A => CO0) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b0)
    (A => CO0) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b1)
    (A => CO0) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b0)
    (A => CO0) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b1)
    (A => CO0) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b0)
    (A => CO0) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b1)
    (A => CO0) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b0)
    (A => CO0) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b1)
    (B => CO0) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b0)
    (B => CO0) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b1)
    (B => CO0) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b0)
    (B => CO0) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b1)
    (B => CO0) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b0)
    (B => CO0) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b1)
    (B => CO0) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b0)
    (B => CO0) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN1 == 1'b1 && CS == 1'b1)
    (CIN0 => CO0) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN1 == 1'b0 && CS == 1'b1)
    (CIN0 => CO0) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN1 == 1'b1 && CS == 1'b1)
    (CIN0 => CO0) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN1 == 1'b0 && CS == 1'b1)
    (CIN0 => CO0) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN1 == 1'b1 && CS == 1'b0)
    (CIN0 => CO0) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN1 == 1'b0 && CS == 1'b0)
    (CIN0 => CO0) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN1 == 1'b1 && CS == 1'b0)
    (CIN0 => CO0) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN1 == 1'b0 && CS == 1'b0)
    (CIN0 => CO0) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b1)
    (A => CO1) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b0)
    (A => CO1) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b1)
    (A => CO1) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b0)
    (A => CO1) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b1)
    (A => CO1) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b0)
    (A => CO1) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b1)
    (A => CO1) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b0)
    (A => CO1) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b1)
    (B => CO1) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b0)
    (B => CO1) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b1)
    (B => CO1) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b0)
    (B => CO1) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b1)
    (B => CO1) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b0)
    (B => CO1) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b1)
    (B => CO1) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b0)
    (B => CO1) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN0 == 1'b1 && CS == 1'b1)
    (CIN1 => CO1) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN0 == 1'b0 && CS == 1'b1)
    (CIN1 => CO1) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN0 == 1'b1 && CS == 1'b1)
    (CIN1 => CO1) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN0 == 1'b0 && CS == 1'b1)
    (CIN1 => CO1) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN0 == 1'b1 && CS == 1'b0)
    (CIN1 => CO1) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN0 == 1'b0 && CS == 1'b0)
    (CIN1 => CO1) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN0 == 1'b1 && CS == 1'b0)
    (CIN1 => CO1) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN0 == 1'b0 && CS == 1'b0)
    (CIN1 => CO1) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN1 == 1'b1 && CS == 1'b0)
    (CIN0 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN1 == 1'b0 && CS == 1'b0)
    (CIN0 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN1 == 1'b1 && CS == 1'b0)
    (CIN0 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN1 == 1'b0 && CS == 1'b0)
    (CIN0 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIN1 == 1'b1 && CS == 1'b0)
    (CIN0 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIN1 == 1'b0 && CS == 1'b0)
    (CIN0 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIN1 == 1'b1 && CS == 1'b0)
    (CIN0 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIN1 == 1'b0 && CS == 1'b0)
    (CIN0 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN0 == 1'b1 && CS == 1'b1)
    (CIN1 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN0 == 1'b0 && CS == 1'b1)
    (CIN1 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN0 == 1'b1 && CS == 1'b1)
    (CIN1 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN0 == 1'b0 && CS == 1'b1)
    (CIN1 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIN0 == 1'b1 && CS == 1'b1)
    (CIN1 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIN0 == 1'b0 && CS == 1'b1)
    (CIN1 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIN0 == 1'b1 && CS == 1'b1)
    (CIN1 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIN0 == 1'b0 && CS == 1'b1)
    (CIN1 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b0)
    (CS => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b0)
    (CS => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b1)
    (CS => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b1)
    (CS => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b1)
    (CS => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b1)
    (CS => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b0)
    (CS => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b0)
    (CS => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FCSICOND1 (A, B, CI0, CI1, CS, S, CON0, CON1);
    input A, B, CI0, CI1, CS;
    output S, CON0, CON1;
    tsmc_mux (I0_out, CI0, CI1, CS);
    xor (I1_out, I0_out, A);
    xor (S, I1_out, B);
    and (I3_out, A, B);
    and (I4_out, B, CI0);
    and (I6_out, CI0, A);
    or (I7_out, I3_out, I4_out, I6_out);
    not (CON0, I7_out);
    and (I9_out, A, B);
    and (I10_out, B, CI1);
    and (I12_out, CI1, A);
    or (I13_out, I9_out, I10_out, I12_out);
    not (CON1, I13_out);

  specify
    if (B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b1)
    (A => CON0) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b0)
    (A => CON0) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b1)
    (A => CON0) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b0)
    (A => CON0) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b1)
    (A => CON0) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b0)
    (A => CON0) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b1)
    (A => CON0) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b0)
    (A => CON0) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b1)
    (B => CON0) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b0)
    (B => CON0) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b1)
    (B => CON0) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b0)
    (B => CON0) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b1)
    (B => CON0) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b0)
    (B => CON0) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b1)
    (B => CON0) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b0)
    (B => CON0) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI1 == 1'b1 && CS == 1'b1)
    (CI0 => CON0) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI1 == 1'b0 && CS == 1'b1)
    (CI0 => CON0) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI1 == 1'b1 && CS == 1'b1)
    (CI0 => CON0) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI1 == 1'b0 && CS == 1'b1)
    (CI0 => CON0) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI1 == 1'b1 && CS == 1'b0)
    (CI0 => CON0) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI1 == 1'b0 && CS == 1'b0)
    (CI0 => CON0) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI1 == 1'b1 && CS == 1'b0)
    (CI0 => CON0) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI1 == 1'b0 && CS == 1'b0)
    (CI0 => CON0) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b1)
    (A => CON1) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b0)
    (A => CON1) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b1)
    (A => CON1) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b0)
    (A => CON1) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b1)
    (A => CON1) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b0)
    (A => CON1) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b1)
    (A => CON1) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b0)
    (A => CON1) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b1)
    (B => CON1) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b0)
    (B => CON1) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b1)
    (B => CON1) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b0)
    (B => CON1) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b1)
    (B => CON1) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b0)
    (B => CON1) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b1)
    (B => CON1) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b0)
    (B => CON1) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI0 == 1'b1 && CS == 1'b1)
    (CI1 => CON1) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI0 == 1'b0 && CS == 1'b1)
    (CI1 => CON1) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI0 == 1'b1 && CS == 1'b1)
    (CI1 => CON1) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI0 == 1'b0 && CS == 1'b1)
    (CI1 => CON1) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI0 == 1'b1 && CS == 1'b0)
    (CI1 => CON1) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI0 == 1'b0 && CS == 1'b0)
    (CI1 => CON1) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI0 == 1'b1 && CS == 1'b0)
    (CI1 => CON1) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI0 == 1'b0 && CS == 1'b0)
    (CI1 => CON1) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CI1 == 1'b1 && CS == 1'b0)
    (CI0 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CI1 == 1'b0 && CS == 1'b0)
    (CI0 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CI1 == 1'b1 && CS == 1'b0)
    (CI0 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CI1 == 1'b0 && CS == 1'b0)
    (CI0 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI1 == 1'b1 && CS == 1'b0)
    (CI0 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI1 == 1'b0 && CS == 1'b0)
    (CI0 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI1 == 1'b1 && CS == 1'b0)
    (CI0 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI1 == 1'b0 && CS == 1'b0)
    (CI0 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CI0 == 1'b1 && CS == 1'b1)
    (CI1 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CI0 == 1'b0 && CS == 1'b1)
    (CI1 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CI0 == 1'b1 && CS == 1'b1)
    (CI1 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CI0 == 1'b0 && CS == 1'b1)
    (CI1 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI0 == 1'b1 && CS == 1'b1)
    (CI1 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI0 == 1'b0 && CS == 1'b1)
    (CI1 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI0 == 1'b1 && CS == 1'b1)
    (CI1 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI0 == 1'b0 && CS == 1'b1)
    (CI1 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1)
    (CS => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1)
    (CS => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0)
    (CS => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0)
    (CS => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0)
    (CS => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0)
    (CS => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1)
    (CS => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1)
    (CS => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FCSICOND2 (A, B, CI0, CI1, CS, S, CON0, CON1);
    input A, B, CI0, CI1, CS;
    output S, CON0, CON1;
    tsmc_mux (I0_out, CI0, CI1, CS);
    xor (I1_out, I0_out, A);
    xor (S, I1_out, B);
    and (I3_out, A, B);
    and (I4_out, B, CI0);
    and (I6_out, CI0, A);
    or (I7_out, I3_out, I4_out, I6_out);
    not (CON0, I7_out);
    and (I9_out, A, B);
    and (I10_out, B, CI1);
    and (I12_out, CI1, A);
    or (I13_out, I9_out, I10_out, I12_out);
    not (CON1, I13_out);

  specify
    if (B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b1)
    (A => CON0) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b0)
    (A => CON0) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b1)
    (A => CON0) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b0)
    (A => CON0) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b1)
    (A => CON0) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b0)
    (A => CON0) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b1)
    (A => CON0) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b0)
    (A => CON0) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b1)
    (B => CON0) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b0)
    (B => CON0) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b1)
    (B => CON0) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b0)
    (B => CON0) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b1)
    (B => CON0) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b0)
    (B => CON0) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b1)
    (B => CON0) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b0)
    (B => CON0) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI1 == 1'b1 && CS == 1'b1)
    (CI0 => CON0) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI1 == 1'b0 && CS == 1'b1)
    (CI0 => CON0) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI1 == 1'b1 && CS == 1'b1)
    (CI0 => CON0) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI1 == 1'b0 && CS == 1'b1)
    (CI0 => CON0) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI1 == 1'b1 && CS == 1'b0)
    (CI0 => CON0) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI1 == 1'b0 && CS == 1'b0)
    (CI0 => CON0) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI1 == 1'b1 && CS == 1'b0)
    (CI0 => CON0) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI1 == 1'b0 && CS == 1'b0)
    (CI0 => CON0) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b1)
    (A => CON1) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b0)
    (A => CON1) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b1)
    (A => CON1) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b0)
    (A => CON1) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b1)
    (A => CON1) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b0)
    (A => CON1) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b1)
    (A => CON1) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b0)
    (A => CON1) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b1)
    (B => CON1) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b0)
    (B => CON1) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b1)
    (B => CON1) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b0)
    (B => CON1) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b1)
    (B => CON1) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b0)
    (B => CON1) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b1)
    (B => CON1) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b0)
    (B => CON1) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI0 == 1'b1 && CS == 1'b1)
    (CI1 => CON1) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI0 == 1'b0 && CS == 1'b1)
    (CI1 => CON1) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI0 == 1'b1 && CS == 1'b1)
    (CI1 => CON1) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI0 == 1'b0 && CS == 1'b1)
    (CI1 => CON1) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI0 == 1'b1 && CS == 1'b0)
    (CI1 => CON1) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI0 == 1'b0 && CS == 1'b0)
    (CI1 => CON1) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI0 == 1'b1 && CS == 1'b0)
    (CI1 => CON1) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI0 == 1'b0 && CS == 1'b0)
    (CI1 => CON1) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CI1 == 1'b1 && CS == 1'b0)
    (CI0 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CI1 == 1'b0 && CS == 1'b0)
    (CI0 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CI1 == 1'b1 && CS == 1'b0)
    (CI0 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CI1 == 1'b0 && CS == 1'b0)
    (CI0 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI1 == 1'b1 && CS == 1'b0)
    (CI0 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI1 == 1'b0 && CS == 1'b0)
    (CI0 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI1 == 1'b1 && CS == 1'b0)
    (CI0 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI1 == 1'b0 && CS == 1'b0)
    (CI0 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CI0 == 1'b1 && CS == 1'b1)
    (CI1 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CI0 == 1'b0 && CS == 1'b1)
    (CI1 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CI0 == 1'b1 && CS == 1'b1)
    (CI1 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CI0 == 1'b0 && CS == 1'b1)
    (CI1 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI0 == 1'b1 && CS == 1'b1)
    (CI1 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI0 == 1'b0 && CS == 1'b1)
    (CI1 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI0 == 1'b1 && CS == 1'b1)
    (CI1 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI0 == 1'b0 && CS == 1'b1)
    (CI1 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1)
    (CS => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1)
    (CS => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0)
    (CS => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0)
    (CS => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0)
    (CS => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0)
    (CS => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1)
    (CS => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1)
    (CS => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FICIND1 (A, B, CIN, S, CO);
    input A, B, CIN;
    output S, CO;
    xor (I0_out, A, B);
    xor (I1_out, I0_out, CIN);
    not (S, I1_out);
    not (I3_out, B);
    not (I4_out, A);
    and (I5_out, I3_out, I4_out);
    not (I6_out, A);
    and (I7_out, I6_out, CIN);
    not (I9_out, B);
    and (I10_out, CIN, I9_out);
    or (I11_out, I5_out, I7_out, I10_out);
    not (CO, I11_out);

  specify
    if (B == 1'b1 && CIN == 1'b1)
    (A => CO) = (0, 0);
    if (B == 1'b0 && CIN == 1'b0)
    (A => CO) = (0, 0);
    if (A == 1'b1 && CIN == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b0 && CIN == 1'b0)
    (B => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CIN => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CIN => CO) = (0, 0);
    if (B == 1'b1 && CIN == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CIN == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CIN == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CIN == 1'b0)
    (A => S) = (0, 0);
    if (A == 1'b1 && CIN == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CIN == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CIN == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CIN == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CIN => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CIN => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1)
    (CIN => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0)
    (CIN => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FICIND2 (A, B, CIN, S, CO);
    input A, B, CIN;
    output S, CO;
    xor (I0_out, A, B);
    xor (I1_out, I0_out, CIN);
    not (S, I1_out);
    not (I3_out, B);
    not (I4_out, A);
    and (I5_out, I3_out, I4_out);
    not (I6_out, A);
    and (I7_out, I6_out, CIN);
    not (I9_out, B);
    and (I10_out, CIN, I9_out);
    or (I11_out, I5_out, I7_out, I10_out);
    not (CO, I11_out);

  specify
    if (B == 1'b1 && CIN == 1'b1)
    (A => CO) = (0, 0);
    if (B == 1'b0 && CIN == 1'b0)
    (A => CO) = (0, 0);
    if (A == 1'b1 && CIN == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b0 && CIN == 1'b0)
    (B => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CIN => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CIN => CO) = (0, 0);
    if (B == 1'b1 && CIN == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CIN == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CIN == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CIN == 1'b0)
    (A => S) = (0, 0);
    if (A == 1'b1 && CIN == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CIN == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CIN == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CIN == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CIN => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CIN => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1)
    (CIN => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0)
    (CIN => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FICOND1 (A, B, CI, S, CON);
    input A, B, CI;
    output S, CON;
    xor (I0_out, A, B);
    xor (S, I0_out, CI);
    and (I2_out, A, B);
    and (I3_out, B, CI);
    and (I5_out, CI, A);
    or (I6_out, I2_out, I3_out, I5_out);
    not (CON, I6_out);

  specify
    if (B == 1'b1 && CI == 1'b0)
    (A => CON) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => CON) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => CON) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => CON) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => CON) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => CON) = (0, 0);
    if (B == 1'b1 && CI == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1)
    (CI => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FICOND2 (A, B, CI, S, CON);
    input A, B, CI;
    output S, CON;
    xor (I0_out, A, B);
    xor (S, I0_out, CI);
    and (I2_out, A, B);
    and (I3_out, B, CI);
    and (I5_out, CI, A);
    or (I6_out, I2_out, I3_out, I5_out);
    not (CON, I6_out);

  specify
    if (B == 1'b1 && CI == 1'b0)
    (A => CON) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => CON) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => CON) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => CON) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => CON) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => CON) = (0, 0);
    if (B == 1'b1 && CI == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1)
    (CI => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FIICOND1 (A, B, C, S, CON0, CON1);
    input A, B, C;
    output S;
    output CON0, CON1;
    xor (I0_out, A, B);
    xor (S, I0_out, C);
    and (I2_out, A, B);
    not (CON0, I2_out);
    or (I4_out, A, B);
    not (CON1, I4_out);

  specify
    if (B == 1'b1 && C == 1'b1)
    (A => CON0) = (0, 0);
    if (B == 1'b1 && C == 1'b0)
    (A => CON0) = (0, 0);
    if (A == 1'b1 && C == 1'b1)
    (B => CON0) = (0, 0);
    if (A == 1'b1 && C == 1'b0)
    (B => CON0) = (0, 0);
    if (B == 1'b0 && C == 1'b1)
    (A => CON1) = (0, 0);
    if (B == 1'b0 && C == 1'b0)
    (A => CON1) = (0, 0);
    if (A == 1'b0 && C == 1'b1)
    (B => CON1) = (0, 0);
    if (A == 1'b0 && C == 1'b0)
    (B => CON1) = (0, 0);
    if (B == 1'b1 && C == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && C == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && C == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && C == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b1 && C == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && C == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && C == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && C == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (C => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FIICOND2 (A, B, C, S, CON0, CON1);
    input A, B, C;
    output S;
    output CON0, CON1;
    xor (I0_out, A, B);
    xor (S, I0_out, C);
    and (I2_out, A, B);
    not (CON0, I2_out);
    or (I4_out, A, B);
    not (CON1, I4_out);

  specify
    if (B == 1'b1 && C == 1'b1)
    (A => CON0) = (0, 0);
    if (B == 1'b1 && C == 1'b0)
    (A => CON0) = (0, 0);
    if (A == 1'b1 && C == 1'b1)
    (B => CON0) = (0, 0);
    if (A == 1'b1 && C == 1'b0)
    (B => CON0) = (0, 0);
    if (B == 1'b0 && C == 1'b1)
    (A => CON1) = (0, 0);
    if (B == 1'b0 && C == 1'b0)
    (A => CON1) = (0, 0);
    if (A == 1'b0 && C == 1'b1)
    (B => CON1) = (0, 0);
    if (A == 1'b0 && C == 1'b0)
    (B => CON1) = (0, 0);
    if (B == 1'b1 && C == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && C == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && C == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && C == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b1 && C == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && C == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && C == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && C == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (C => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GAN2D1 (A1, A2, Z);
    input A1, A2;
    output Z;
    and (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GAN2D2 (A1, A2, Z);
    input A1, A2;
    output Z;
    and (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GAOI22D1 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GBUFFD1 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GBUFFD2 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GBUFFD3 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GBUFFD4 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GBUFFD8 (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GDCAP;
    // No function
endmodule
`endcelldefine

`celldefine
module GDCAP10;
    // No function
endmodule
`endcelldefine

`celldefine
module GDFQD1 (D, CP, Q);
    input D, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
  `endif

    not (nD, D);

  // Timing logics defined for default constraint check
  pullup  (CP_check);
  pullup  (D_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:D)) = (0, 0);
    $width (posedge CP &&& D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module GINVD1 (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GINVD2 (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GINVD3 (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GINVD4 (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GINVD8 (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GMUX2D1 (I0, I1, S, Z);
    input I0, I1, S;
    output Z;
    tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GMUX2D2 (I0, I1, S, Z);
    input I0, I1, S;
    output Z;
    tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GND2D1 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GND2D2 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GND2D3 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GND2D4 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GND3D1 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    and (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GND3D2 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    and (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GNR2D1 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    or (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GNR2D2 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    or (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GOR2D1 (A1, A2, Z);
    input A1, A2;
    output Z;
    or (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GOR2D2 (A1, A2, Z);
    input A1, A2;
    output Z;
    or (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GXNR2D1 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    xor (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    if (A2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0)
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GXNR2D2 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    xor (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    if (A2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0)
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GXOR2D1 (A1, A2, Z);
    input A1, A2;
    output Z;
    xor (Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GXOR2D2 (A1, A2, Z);
    input A1, A2;
    output Z;
    xor (Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module HA1D0 (A, B, S, CO);
    input A, B;
    output S, CO;
    xor (S, A, B);
    and (CO, A, B);

  specify
    (A => CO) = (0, 0);
    (B => CO) = (0, 0);
    if (B == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1)
    (B => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module HA1D1 (A, B, S, CO);
    input A, B;
    output S, CO;
    xor (S, A, B);
    and (CO, A, B);

  specify
    (A => CO) = (0, 0);
    (B => CO) = (0, 0);
    if (B == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1)
    (B => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module HA1D2 (A, B, S, CO);
    input A, B;
    output S, CO;
    xor (S, A, B);
    and (CO, A, B);

  specify
    (A => CO) = (0, 0);
    (B => CO) = (0, 0);
    if (B == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1)
    (B => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module HA1D4 (A, B, S, CO);
    input A, B;
    output S, CO;
    xor (S, A, B);
    and (CO, A, B);

  specify
    (A => CO) = (0, 0);
    (B => CO) = (0, 0);
    if (B == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1)
    (B => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module HCOSCIND1 (A, CIN, CS, S, CO);
    input A, CIN, CS;
    output S, CO;
    xor (I0_out, A, CIN);
    not (I1_out, I0_out);
    tsmc_mux (S, A, I1_out, CS);
    not (I2_out, CIN);
    and (CO, I2_out, A);

  specify
    if (CIN == 1'b0 && CS == 1'b1)
    (A => CO) = (0, 0);
    if (CIN == 1'b0 && CS == 1'b0)
    (A => CO) = (0, 0);
    if (A == 1'b1 && CS == 1'b1)
    (CIN => CO) = (0, 0);
    if (A == 1'b1 && CS == 1'b0)
    (CIN => CO) = (0, 0);
    if (CIN == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (CIN == 1'b1 && CS == 1'b0)
    (A => S) = (0, 0);
    if (CIN == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (CIN == 1'b0 && CS == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b1 && CS == 1'b1)
    (CIN => S) = (0, 0);
    if (A == 1'b0 && CS == 1'b1)
    (CIN => S) = (0, 0);
    if (A == 1'b0 && CIN == 1'b0)
    (CS => S) = (0, 0);
    if (A == 1'b1 && CIN == 1'b0)
    (CS => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module HCOSCIND2 (A, CIN, CS, S, CO);
    input A, CIN, CS;
    output S, CO;
    xor (I0_out, A, CIN);
    not (I1_out, I0_out);
    tsmc_mux (S, A, I1_out, CS);
    not (I2_out, CIN);
    and (CO, I2_out, A);

  specify
    if (CIN == 1'b0 && CS == 1'b1)
    (A => CO) = (0, 0);
    if (CIN == 1'b0 && CS == 1'b0)
    (A => CO) = (0, 0);
    if (A == 1'b1 && CS == 1'b1)
    (CIN => CO) = (0, 0);
    if (A == 1'b1 && CS == 1'b0)
    (CIN => CO) = (0, 0);
    if (CIN == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (CIN == 1'b1 && CS == 1'b0)
    (A => S) = (0, 0);
    if (CIN == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (CIN == 1'b0 && CS == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b1 && CS == 1'b1)
    (CIN => S) = (0, 0);
    if (A == 1'b0 && CS == 1'b1)
    (CIN => S) = (0, 0);
    if (A == 1'b0 && CIN == 1'b0)
    (CS => S) = (0, 0);
    if (A == 1'b1 && CIN == 1'b0)
    (CS => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module HCOSCOND1 (A, CI, CS, S, CON);
    input A, CI, CS;
    output S, CON;
    xor (I0_out, A, CI);
    tsmc_mux (S, A, I0_out, CS);
    and (I1_out, A, CI);
    not (CON, I1_out);

  specify
    if (CI == 1'b1 && CS == 1'b1)
    (A => CON) = (0, 0);
    if (CI == 1'b1 && CS == 1'b0)
    (A => CON) = (0, 0);
    if (A == 1'b1 && CS == 1'b1)
    (CI => CON) = (0, 0);
    if (A == 1'b1 && CS == 1'b0)
    (CI => CON) = (0, 0);
    if (CI == 1'b1 && CS == 1'b0)
    (A => S) = (0, 0);
    if (CI == 1'b0 && CS == 1'b1)
    (A => S) = (0, 0);
    if (CI == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (CI == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b0 && CS == 1'b1)
    (CI => S) = (0, 0);
    if (A == 1'b1 && CS == 1'b1)
    (CI => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (CS => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b1)
    (CS => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module HCOSCOND2 (A, CI, CS, S, CON);
    input A, CI, CS;
    output S, CON;
    xor (I0_out, A, CI);
    tsmc_mux (S, A, I0_out, CS);
    and (I1_out, A, CI);
    not (CON, I1_out);

  specify
    if (CI == 1'b1 && CS == 1'b1)
    (A => CON) = (0, 0);
    if (CI == 1'b1 && CS == 1'b0)
    (A => CON) = (0, 0);
    if (A == 1'b1 && CS == 1'b1)
    (CI => CON) = (0, 0);
    if (A == 1'b1 && CS == 1'b0)
    (CI => CON) = (0, 0);
    if (CI == 1'b1 && CS == 1'b0)
    (A => S) = (0, 0);
    if (CI == 1'b0 && CS == 1'b1)
    (A => S) = (0, 0);
    if (CI == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (CI == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b0 && CS == 1'b1)
    (CI => S) = (0, 0);
    if (A == 1'b1 && CS == 1'b1)
    (CI => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (CS => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b1)
    (CS => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module HICIND1 (A, CIN, S, CO);
    input A, CIN;
    output S, CO;
    xor (I0_out, A, CIN);
    not (S, I0_out);
    not (I1_out, CIN);
    and (CO, I1_out, A);

  specify
    (A => CO) = (0, 0);
    (CIN => CO) = (0, 0);
    if (CIN == 1'b1)
    (A => S) = (0, 0);
    if (CIN == 1'b0)
    (A => S) = (0, 0);
    if (A == 1'b1)
    (CIN => S) = (0, 0);
    if (A == 1'b0)
    (CIN => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module HICIND2 (A, CIN, S, CO);
    input A, CIN;
    output S, CO;
    xor (I0_out, A, CIN);
    not (S, I0_out);
    not (I1_out, CIN);
    and (CO, I1_out, A);

  specify
    (A => CO) = (0, 0);
    (CIN => CO) = (0, 0);
    if (CIN == 1'b1)
    (A => S) = (0, 0);
    if (CIN == 1'b0)
    (A => S) = (0, 0);
    if (A == 1'b1)
    (CIN => S) = (0, 0);
    if (A == 1'b0)
    (CIN => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module HICOND1 (A, CI, S, CON);
    input A, CI;
    output S, CON;
    xor (S, A, CI);
    and (I1_out, A, CI);
    not (CON, I1_out);

  specify
    (A => CON) = (0, 0);
    (CI => CON) = (0, 0);
    if (CI == 1'b0)
    (A => S) = (0, 0);
    if (CI == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b1)
    (CI => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module HICOND2 (A, CI, S, CON);
    input A, CI;
    output S, CON;
    xor (S, A, CI);
    and (I1_out, A, CI);
    not (CON, I1_out);

  specify
    (A => CON) = (0, 0);
    (CI => CON) = (0, 0);
    if (CI == 1'b0)
    (A => S) = (0, 0);
    if (CI == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b1)
    (CI => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IAO21D0 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    not (I0_out, A1);
    not (I1_out, A2);
    and (I2_out, I1_out, I0_out);
    or (Z, I2_out, B);
    not (ZN, Z);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IAO21D1 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    not (I0_out, A1);
    not (I1_out, A2);
    and (I2_out, I1_out, I0_out);
    or (Z, I2_out, B);
    not (ZN, Z);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IAO21D2 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    not (I0_out, A1);
    not (I1_out, A2);
    and (I2_out, I1_out, I0_out);
    or (Z, I2_out, B);
    not (ZN, Z);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IAO21D4 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    not (I0_out, A1);
    not (I1_out, A2);
    and (I2_out, I1_out, I0_out);
    or (Z, I2_out, B);
    not (ZN, Z);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IAO22D0 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    not (I0_out, A1);
    not (I1_out, A2);
    and (I2_out, I1_out, I0_out);
    and (I3_out, B1, B2);
    or (I4_out, I3_out, I2_out);
    not (ZN, I4_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IAO22D1 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    not (I0_out, A1);
    not (I1_out, A2);
    and (I2_out, I1_out, I0_out);
    and (I3_out, B1, B2);
    or (I4_out, I3_out, I2_out);
    not (ZN, I4_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IAO22D2 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    not (I0_out, A1);
    not (I1_out, A2);
    and (I2_out, I1_out, I0_out);
    and (I3_out, B1, B2);
    or (I4_out, I3_out, I2_out);
    not (ZN, I4_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IAO22D4 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    not (I0_out, A1);
    not (I1_out, A2);
    and (I2_out, I1_out, I0_out);
    and (I3_out, B1, B2);
    or (I4_out, I3_out, I2_out);
    not (ZN, I4_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IIND4D0 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    not (I0_out, A1);
    not (I1_out, A2);
    and (I2_out, I0_out, I1_out, B1, B2);
    not (ZN, I2_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IIND4D1 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    not (I0_out, A1);
    not (I1_out, A2);
    and (I2_out, I0_out, I1_out, B1, B2);
    not (ZN, I2_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IIND4D2 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    not (I0_out, A1);
    not (I1_out, A2);
    and (I2_out, I0_out, I1_out, B1, B2);
    not (ZN, I2_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IIND4D4 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    not (I0_out, A1);
    not (I1_out, A2);
    and (I2_out, I0_out, I1_out, B1, B2);
    not (ZN, I2_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IINR4D0 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    not (I0_out, A1);
    not (I1_out, A2);
    or (I2_out, I0_out, I1_out, B1, B2);
    not (ZN, I2_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IINR4D1 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    not (I0_out, A1);
    not (I1_out, A2);
    or (I2_out, I0_out, I1_out, B1, B2);
    not (ZN, I2_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IINR4D2 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    not (I0_out, A1);
    not (I1_out, A2);
    or (I2_out, I0_out, I1_out, B1, B2);
    not (ZN, I2_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IINR4D4 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    not (I0_out, A1);
    not (I1_out, A2);
    or (I2_out, I0_out, I1_out, B1, B2);
    not (ZN, I2_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND2D0 (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not (I0_out, A1);
    and (I1_out, I0_out, B1);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND2D1 (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not (I0_out, A1);
    and (I1_out, I0_out, B1);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND2D2 (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not (I0_out, A1);
    and (I1_out, I0_out, B1);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND2D4 (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not (I0_out, A1);
    and (I1_out, I0_out, B1);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND3D0 (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
    not (I0_out, A1);
    and (I1_out, I0_out, B1, B2);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND3D1 (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
    not (I0_out, A1);
    and (I1_out, I0_out, B1, B2);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND3D2 (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
    not (I0_out, A1);
    and (I1_out, I0_out, B1, B2);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND3D4 (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
    not (I0_out, A1);
    and (I1_out, I0_out, B1, B2);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND4D0 (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
    not (I0_out, A1);
    and (I1_out, I0_out, B1, B2, B3);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND4D1 (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
    not (I0_out, A1);
    and (I1_out, I0_out, B1, B2, B3);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND4D2 (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
    not (I0_out, A1);
    and (I1_out, I0_out, B1, B2, B3);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND4D4 (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
    not (I0_out, A1);
    and (I1_out, I0_out, B1, B2, B3);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR2D0 (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not (I0_out, A1);
    or (I1_out, I0_out, B1);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR2D1 (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not (I0_out, A1);
    or (I1_out, I0_out, B1);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR2D2 (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not (I0_out, A1);
    or (I1_out, I0_out, B1);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR2D4 (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not (I0_out, A1);
    or (I1_out, I0_out, B1);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR2XD0 (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not (I0_out, A1);
    or (I1_out, I0_out, B1);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR2XD1 (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not (I0_out, A1);
    or (I1_out, I0_out, B1);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR2XD2 (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not (I0_out, A1);
    or (I1_out, I0_out, B1);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR2XD4 (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not (I0_out, A1);
    or (I1_out, I0_out, B1);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR3D0 (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
    not (I0_out, A1);
    or (I1_out, I0_out, B1, B2);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR3D1 (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
    not (I0_out, A1);
    or (I1_out, I0_out, B1, B2);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR3D2 (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
    not (I0_out, A1);
    or (I1_out, I0_out, B1, B2);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR3D4 (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
    not (I0_out, A1);
    or (I1_out, I0_out, B1, B2);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR4D0 (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
    not (I0_out, A1);
    or (I1_out, I0_out, B1, B2, B3);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR4D1 (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
    not (I0_out, A1);
    or (I1_out, I0_out, B1, B2, B3);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR4D2 (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
    not (I0_out, A1);
    or (I1_out, I0_out, B1, B2, B3);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR4D4 (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
    not (I0_out, A1);
    or (I1_out, I0_out, B1, B2, B3);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INVD0 (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INVD1 (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INVD12 (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INVD16 (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INVD2 (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INVD20 (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INVD24 (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INVD3 (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INVD4 (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INVD6 (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INVD8 (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IOA21D0 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    and (I0_out, A1, A2);
    not (I1_out, I0_out);
    and (I2_out, I1_out, B);
    not (ZN, I2_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IOA21D1 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    and (I0_out, A1, A2);
    not (I1_out, I0_out);
    and (I2_out, I1_out, B);
    not (ZN, I2_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IOA21D2 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    and (I0_out, A1, A2);
    not (I1_out, I0_out);
    and (I2_out, I1_out, B);
    not (ZN, I2_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IOA21D4 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    and (I0_out, A1, A2);
    not (I1_out, I0_out);
    and (I2_out, I1_out, B);
    not (ZN, I2_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IOA22D0 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or (I0_out, B1, B2);
    not (I1_out, I0_out);
    and (I2_out, A1, A2);
    or (ZN, I1_out, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IOA22D1 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or (I0_out, B1, B2);
    not (I1_out, I0_out);
    and (I2_out, A1, A2);
    or (ZN, I1_out, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IOA22D2 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or (I0_out, B1, B2);
    not (I1_out, I0_out);
    and (I2_out, A1, A2);
    or (ZN, I1_out, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IOA22D4 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or (I0_out, B1, B2);
    not (I1_out, I0_out);
    and (I2_out, A1, A2);
    or (ZN, I1_out, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LHCND1 (D, E, CDN, Q, QN);
    input D, E, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, E_d;
        pullup (SDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nE, E);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (D == 1'b1 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    if (D == 1'b1 && E == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    $width (negedge CDN &&& D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_nE_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0,0, notifier, , , CDN_d, E_d);
    `else
      $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0, notifier);
      $hold (negedge E &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0, notifier);
    $hold (negedge E &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCND2 (D, E, CDN, Q, QN);
    input D, E, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, E_d;
        pullup (SDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nE, E);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (D == 1'b1 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    if (D == 1'b1 && E == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    $width (negedge CDN &&& D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_nE_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0,0, notifier, , , CDN_d, E_d);
    `else
      $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0, notifier);
      $hold (negedge E &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0, notifier);
    $hold (negedge E &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCND4 (D, E, CDN, Q, QN);
    input D, E, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, E_d;
        pullup (SDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nE, E);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (D == 1'b1 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    if (D == 1'b1 && E == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    $width (negedge CDN &&& D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_nE_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0,0, notifier, , , CDN_d, E_d);
    `else
      $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0, notifier);
      $hold (negedge E &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0, notifier);
    $hold (negedge E &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCNQD1 (D, E, CDN, Q);
    input D, E, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, E_d;
        pullup (SDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nE, E);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (D == 1'b1 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    $width (negedge CDN &&& D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_nE_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0,0, notifier, , , CDN_d, E_d);
    `else
      $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0, notifier);
      $hold (negedge E &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0, notifier);
    $hold (negedge E &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCNQD2 (D, E, CDN, Q);
    input D, E, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, E_d;
        pullup (SDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nE, E);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (D == 1'b1 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    $width (negedge CDN &&& D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_nE_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0,0, notifier, , , CDN_d, E_d);
    `else
      $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0, notifier);
      $hold (negedge E &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0, notifier);
    $hold (negedge E &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCNQD4 (D, E, CDN, Q);
    input D, E, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, E_d;
        pullup (SDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nE, E);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (D == 1'b1 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    $width (negedge CDN &&& D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_nE_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0,0, notifier, , , CDN_d, E_d);
    `else
      $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0, notifier);
      $hold (negedge E &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0, notifier);
    $hold (negedge E &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCSND1 (D, E, CDN, SDN, Q, QN);
    input D, E, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, E_d;
        tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_nE_SDN_SDFCHK, D_nE_SDN, 1'b1);
    tsmc_xbuf (nD_nE_SDN_SDFCHK, nD_nE_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_nE_SDFCHK, CDN_D_nE, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SDFCHK, CDN_nD_nE, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nE, E);
    and (D_nE_SDN, D, nE, SDN);
    and (nD_nE_SDN, nD, nE, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_D_nE, CDN, D, nE);
    and (CDN_nD_nE, CDN, nD, nE);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (D == 1'b1 && E == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b1 && E == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && E == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge CDN &&& D_nE_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_nE_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nD_nE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, E_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0, notifier);
      $hold (negedge E &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (negedge E &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0, notifier);
    $hold (negedge E &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (negedge E &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCSND2 (D, E, CDN, SDN, Q, QN);
    input D, E, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, E_d;
        tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_nE_SDN_SDFCHK, D_nE_SDN, 1'b1);
    tsmc_xbuf (nD_nE_SDN_SDFCHK, nD_nE_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_nE_SDFCHK, CDN_D_nE, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SDFCHK, CDN_nD_nE, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nE, E);
    and (D_nE_SDN, D, nE, SDN);
    and (nD_nE_SDN, nD, nE, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_D_nE, CDN, D, nE);
    and (CDN_nD_nE, CDN, nD, nE);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (D == 1'b1 && E == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b1 && E == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && E == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge CDN &&& D_nE_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_nE_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nD_nE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, E_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0, notifier);
      $hold (negedge E &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (negedge E &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0, notifier);
    $hold (negedge E &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (negedge E &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCSND4 (D, E, CDN, SDN, Q, QN);
    input D, E, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, E_d;
        tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_nE_SDN_SDFCHK, D_nE_SDN, 1'b1);
    tsmc_xbuf (nD_nE_SDN_SDFCHK, nD_nE_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_nE_SDFCHK, CDN_D_nE, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SDFCHK, CDN_nD_nE, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nE, E);
    and (D_nE_SDN, D, nE, SDN);
    and (nD_nE_SDN, nD, nE, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_D_nE, CDN, D, nE);
    and (CDN_nD_nE, CDN, nD, nE);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (D == 1'b1 && E == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b1 && E == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && E == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge CDN &&& D_nE_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_nE_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nD_nE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, E_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0, notifier);
      $hold (negedge E &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (negedge E &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0, notifier);
    $hold (negedge E &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (negedge E &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCSNQD1 (D, E, CDN, SDN, Q);
    input D, E, CDN, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, E_d;
        tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_nE_SDN_SDFCHK, D_nE_SDN, 1'b1);
    tsmc_xbuf (nD_nE_SDN_SDFCHK, nD_nE_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_nE_SDFCHK, CDN_D_nE, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SDFCHK, CDN_nD_nE, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nE, E);
    and (D_nE_SDN, D, nE, SDN);
    and (nD_nE_SDN, nD, nE, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_D_nE, CDN, D, nE);
    and (CDN_nD_nE, CDN, nD, nE);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (D == 1'b1 && E == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (negedge CDN &&& D_nE_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_nE_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nD_nE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, E_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0, notifier);
      $hold (negedge E &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (negedge E &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0, notifier);
    $hold (negedge E &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (negedge E &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCSNQD2 (D, E, CDN, SDN, Q);
    input D, E, CDN, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, E_d;
        tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_nE_SDN_SDFCHK, D_nE_SDN, 1'b1);
    tsmc_xbuf (nD_nE_SDN_SDFCHK, nD_nE_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_nE_SDFCHK, CDN_D_nE, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SDFCHK, CDN_nD_nE, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nE, E);
    and (D_nE_SDN, D, nE, SDN);
    and (nD_nE_SDN, nD, nE, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_D_nE, CDN, D, nE);
    and (CDN_nD_nE, CDN, nD, nE);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (D == 1'b1 && E == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (negedge CDN &&& D_nE_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_nE_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nD_nE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, E_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0, notifier);
      $hold (negedge E &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (negedge E &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0, notifier);
    $hold (negedge E &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (negedge E &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCSNQD4 (D, E, CDN, SDN, Q);
    input D, E, CDN, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, E_d;
        tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_nE_SDN_SDFCHK, D_nE_SDN, 1'b1);
    tsmc_xbuf (nD_nE_SDN_SDFCHK, nD_nE_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_nE_SDFCHK, CDN_D_nE, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SDFCHK, CDN_nD_nE, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    not (nE, E);
    and (D_nE_SDN, D, nE, SDN);
    and (nD_nE_SDN, nD, nE, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_D_nE, CDN, D, nE);
    and (CDN_nD_nE, CDN, nD, nE);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (D == 1'b1 && E == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (negedge CDN &&& D_nE_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_nE_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nD_nE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, E_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0, notifier);
      $hold (negedge E &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (negedge E &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0, notifier);
    $hold (negedge E &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (negedge E &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHD1 (D, E, Q, QN);
    input D, E;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, E_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
  `endif

    not (nD, D);

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    $width (posedge E &&& D_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge E, posedge D, 0, 0, notifier,,, E_d, D_d);
    $setuphold (negedge E, negedge D, 0, 0, notifier,,, E_d, D_d);
  `else
    $setuphold (negedge E, posedge D, 0, 0, notifier);
    $setuphold (negedge E, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHD2 (D, E, Q, QN);
    input D, E;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, E_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
  `endif

    not (nD, D);

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    $width (posedge E &&& D_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge E, posedge D, 0, 0, notifier,,, E_d, D_d);
    $setuphold (negedge E, negedge D, 0, 0, notifier,,, E_d, D_d);
  `else
    $setuphold (negedge E, posedge D, 0, 0, notifier);
    $setuphold (negedge E, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHD4 (D, E, Q, QN);
    input D, E;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, E_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
  `endif

    not (nD, D);

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    $width (posedge E &&& D_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge E, posedge D, 0, 0, notifier,,, E_d, D_d);
    $setuphold (negedge E, negedge D, 0, 0, notifier,,, E_d, D_d);
  `else
    $setuphold (negedge E, posedge D, 0, 0, notifier);
    $setuphold (negedge E, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHQD1 (D, E, Q);
    input D, E;
    output Q;
    reg notifier;
    `ifdef NTC
        wire D_d, E_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
  `endif

    not (nD, D);

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    $width (posedge E &&& D_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge E, posedge D, 0, 0, notifier,,, E_d, D_d);
    $setuphold (negedge E, negedge D, 0, 0, notifier,,, E_d, D_d);
  `else
    $setuphold (negedge E, posedge D, 0, 0, notifier);
    $setuphold (negedge E, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHQD2 (D, E, Q);
    input D, E;
    output Q;
    reg notifier;
    `ifdef NTC
        wire D_d, E_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
  `endif

    not (nD, D);

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    $width (posedge E &&& D_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge E, posedge D, 0, 0, notifier,,, E_d, D_d);
    $setuphold (negedge E, negedge D, 0, 0, notifier,,, E_d, D_d);
  `else
    $setuphold (negedge E, posedge D, 0, 0, notifier);
    $setuphold (negedge E, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHQD4 (D, E, Q);
    input D, E;
    output Q;
    reg notifier;
    `ifdef NTC
        wire D_d, E_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
  `endif

    not (nD, D);

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    $width (posedge E &&& D_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge E, posedge D, 0, 0, notifier,,, E_d, D_d);
    $setuphold (negedge E, negedge D, 0, 0, notifier,,, E_d, D_d);
  `else
    $setuphold (negedge E, posedge D, 0, 0, notifier);
    $setuphold (negedge E, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHSND1 (D, E, SDN, Q, QN);
    input D, E, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, E_d;
        pullup (CDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_dla (Q_buf, D, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
  `endif

    not (nD, D);
    not (nE, E);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);

  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge E &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nD_nE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0, notifier);
      $hold (negedge E &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0, notifier);
    $hold (negedge E &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHSND2 (D, E, SDN, Q, QN);
    input D, E, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, E_d;
        pullup (CDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_dla (Q_buf, D, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
  `endif

    not (nD, D);
    not (nE, E);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);

  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge E &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nD_nE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0, notifier);
      $hold (negedge E &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0, notifier);
    $hold (negedge E &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHSND4 (D, E, SDN, Q, QN);
    input D, E, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, E_d;
        pullup (CDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_dla (Q_buf, D, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
  `endif

    not (nD, D);
    not (nE, E);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);

  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge E &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nD_nE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0, notifier);
      $hold (negedge E &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0, notifier);
    $hold (negedge E &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHSNQD1 (D, E, SDN, Q);
    input D, E, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, E_d;
        pullup (CDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_dla (Q_buf, D, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
  `endif

    not (nD, D);
    not (nE, E);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);

  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (posedge E &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nD_nE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0, notifier);
      $hold (negedge E &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0, notifier);
    $hold (negedge E &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHSNQD2 (D, E, SDN, Q);
    input D, E, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, E_d;
        pullup (CDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_dla (Q_buf, D, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
  `endif

    not (nD, D);
    not (nE, E);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);

  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (posedge E &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nD_nE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0, notifier);
      $hold (negedge E &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0, notifier);
    $hold (negedge E &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHSNQD4 (D, E, SDN, Q);
    input D, E, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, E_d;
        pullup (CDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_dla (Q_buf, D, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
  `endif

    not (nD, D);
    not (nE, E);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);

  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (posedge E &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nD_nE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0, notifier);
      $hold (negedge E &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0, notifier);
    $hold (negedge E &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCND1 (D, EN, CDN, Q, QN);
    input D, EN, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, EN_d;
        pullup (SDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (D == 1'b1 && EN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    if (D == 1'b1 && EN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    $width (negedge CDN &&& D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_EN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0,0, notifier, , , CDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0, notifier);
      $hold (posedge EN &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0, notifier);
    $hold (posedge EN &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCND2 (D, EN, CDN, Q, QN);
    input D, EN, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, EN_d;
        pullup (SDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (D == 1'b1 && EN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    if (D == 1'b1 && EN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    $width (negedge CDN &&& D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_EN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0,0, notifier, , , CDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0, notifier);
      $hold (posedge EN &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0, notifier);
    $hold (posedge EN &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCND4 (D, EN, CDN, Q, QN);
    input D, EN, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, EN_d;
        pullup (SDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (D == 1'b1 && EN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    if (D == 1'b1 && EN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    $width (negedge CDN &&& D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_EN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0,0, notifier, , , CDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0, notifier);
      $hold (posedge EN &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0, notifier);
    $hold (posedge EN &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCNQD1 (D, EN, CDN, Q);
    input D, EN, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, EN_d;
        pullup (SDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (D == 1'b1 && EN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    $width (negedge CDN &&& D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_EN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0,0, notifier, , , CDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0, notifier);
      $hold (posedge EN &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0, notifier);
    $hold (posedge EN &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCNQD2 (D, EN, CDN, Q);
    input D, EN, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, EN_d;
        pullup (SDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (D == 1'b1 && EN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    $width (negedge CDN &&& D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_EN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0,0, notifier, , , CDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0, notifier);
      $hold (posedge EN &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0, notifier);
    $hold (posedge EN &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCNQD4 (D, EN, CDN, Q);
    input D, EN, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, EN_d;
        pullup (SDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (D == 1'b1 && EN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    $width (negedge CDN &&& D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_EN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0,0, notifier, , , CDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0, notifier);
      $hold (posedge EN &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0, notifier);
    $hold (posedge EN &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCSND1 (D, EN, CDN, SDN, Q, QN);
    input D, EN, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, EN_d;
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_EN_SDN_SDFCHK, D_EN_SDN, 1'b1);
    tsmc_xbuf (nD_EN_SDN_SDFCHK, nD_EN_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_EN_SDFCHK, CDN_D_EN, 1'b1);
    tsmc_xbuf (CDN_nD_EN_SDFCHK, CDN_nD_EN, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    and (D_EN_SDN, D, EN, SDN);
    and (nD_EN_SDN, nD, EN, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_D_EN, CDN, D, EN);
    and (CDN_nD_EN, CDN, nD, EN);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (D == 1'b1 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b1 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && EN == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge CDN &&& D_EN_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_EN_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nD_EN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, EN_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0, notifier);
      $hold (posedge EN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (posedge EN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0, notifier);
    $hold (posedge EN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (posedge EN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCSND2 (D, EN, CDN, SDN, Q, QN);
    input D, EN, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, EN_d;
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_EN_SDN_SDFCHK, D_EN_SDN, 1'b1);
    tsmc_xbuf (nD_EN_SDN_SDFCHK, nD_EN_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_EN_SDFCHK, CDN_D_EN, 1'b1);
    tsmc_xbuf (CDN_nD_EN_SDFCHK, CDN_nD_EN, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    and (D_EN_SDN, D, EN, SDN);
    and (nD_EN_SDN, nD, EN, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_D_EN, CDN, D, EN);
    and (CDN_nD_EN, CDN, nD, EN);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (D == 1'b1 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b1 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && EN == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge CDN &&& D_EN_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_EN_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nD_EN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, EN_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0, notifier);
      $hold (posedge EN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (posedge EN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0, notifier);
    $hold (posedge EN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (posedge EN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCSND4 (D, EN, CDN, SDN, Q, QN);
    input D, EN, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, EN_d;
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_EN_SDN_SDFCHK, D_EN_SDN, 1'b1);
    tsmc_xbuf (nD_EN_SDN_SDFCHK, nD_EN_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_EN_SDFCHK, CDN_D_EN, 1'b1);
    tsmc_xbuf (CDN_nD_EN_SDFCHK, CDN_nD_EN, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    and (D_EN_SDN, D, EN, SDN);
    and (nD_EN_SDN, nD, EN, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_D_EN, CDN, D, EN);
    and (CDN_nD_EN, CDN, nD, EN);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (D == 1'b1 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b1 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && EN == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge CDN &&& D_EN_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_EN_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nD_EN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, EN_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0, notifier);
      $hold (posedge EN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (posedge EN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0, notifier);
    $hold (posedge EN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (posedge EN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCSNQD1 (D, EN, CDN, SDN, Q);
    input D, EN, CDN, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, EN_d;
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_EN_SDN_SDFCHK, D_EN_SDN, 1'b1);
    tsmc_xbuf (nD_EN_SDN_SDFCHK, nD_EN_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_EN_SDFCHK, CDN_D_EN, 1'b1);
    tsmc_xbuf (CDN_nD_EN_SDFCHK, CDN_nD_EN, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    and (D_EN_SDN, D, EN, SDN);
    and (nD_EN_SDN, nD, EN, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_D_EN, CDN, D, EN);
    and (CDN_nD_EN, CDN, nD, EN);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (D == 1'b1 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (negedge CDN &&& D_EN_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_EN_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nD_EN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, EN_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0, notifier);
      $hold (posedge EN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (posedge EN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0, notifier);
    $hold (posedge EN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (posedge EN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCSNQD2 (D, EN, CDN, SDN, Q);
    input D, EN, CDN, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, EN_d;
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_EN_SDN_SDFCHK, D_EN_SDN, 1'b1);
    tsmc_xbuf (nD_EN_SDN_SDFCHK, nD_EN_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_EN_SDFCHK, CDN_D_EN, 1'b1);
    tsmc_xbuf (CDN_nD_EN_SDFCHK, CDN_nD_EN, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    and (D_EN_SDN, D, EN, SDN);
    and (nD_EN_SDN, nD, EN, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_D_EN, CDN, D, EN);
    and (CDN_nD_EN, CDN, nD, EN);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (D == 1'b1 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (negedge CDN &&& D_EN_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_EN_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nD_EN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, EN_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0, notifier);
      $hold (posedge EN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (posedge EN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0, notifier);
    $hold (posedge EN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (posedge EN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCSNQD4 (D, EN, CDN, SDN, Q);
    input D, EN, CDN, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, EN_d;
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_EN_SDN_SDFCHK, D_EN_SDN, 1'b1);
    tsmc_xbuf (nD_EN_SDN_SDFCHK, nD_EN_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_EN_SDFCHK, CDN_D_EN, 1'b1);
    tsmc_xbuf (CDN_nD_EN_SDFCHK, CDN_nD_EN, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
  `endif

    not (nD, D);
    and (D_EN_SDN, D, EN, SDN);
    and (nD_EN_SDN, nD, EN, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_D_EN, CDN, D, EN);
    and (CDN_nD_EN, CDN, nD, EN);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);

  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (D == 1'b1 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (negedge CDN &&& D_EN_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_EN_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nD_EN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, EN_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0, notifier);
      $hold (posedge EN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (posedge EN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0, notifier);
    $hold (posedge EN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (posedge EN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LND1 (D, EN, Q, QN);
    input D, EN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, EN_d;
        pullup (CDN);
        pullup (SDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
  `endif

    not (nD, D);

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    $width (negedge EN &&& D_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge EN, posedge D, 0, 0, notifier,,, EN_d, D_d);
    $setuphold (posedge EN, negedge D, 0, 0, notifier,,, EN_d, D_d);
  `else
    $setuphold (posedge EN, posedge D, 0, 0, notifier);
    $setuphold (posedge EN, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LND2 (D, EN, Q, QN);
    input D, EN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, EN_d;
        pullup (CDN);
        pullup (SDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
  `endif

    not (nD, D);

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    $width (negedge EN &&& D_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge EN, posedge D, 0, 0, notifier,,, EN_d, D_d);
    $setuphold (posedge EN, negedge D, 0, 0, notifier,,, EN_d, D_d);
  `else
    $setuphold (posedge EN, posedge D, 0, 0, notifier);
    $setuphold (posedge EN, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LND4 (D, EN, Q, QN);
    input D, EN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, EN_d;
        pullup (CDN);
        pullup (SDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
  `endif

    not (nD, D);

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    $width (negedge EN &&& D_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge EN, posedge D, 0, 0, notifier,,, EN_d, D_d);
    $setuphold (posedge EN, negedge D, 0, 0, notifier,,, EN_d, D_d);
  `else
    $setuphold (posedge EN, posedge D, 0, 0, notifier);
    $setuphold (posedge EN, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNQD1 (D, EN, Q);
    input D, EN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire D_d, EN_d;
        pullup (CDN);
        pullup (SDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
  `endif

    not (nD, D);

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    $width (negedge EN &&& D_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge EN, posedge D, 0, 0, notifier,,, EN_d, D_d);
    $setuphold (posedge EN, negedge D, 0, 0, notifier,,, EN_d, D_d);
  `else
    $setuphold (posedge EN, posedge D, 0, 0, notifier);
    $setuphold (posedge EN, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNQD2 (D, EN, Q);
    input D, EN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire D_d, EN_d;
        pullup (CDN);
        pullup (SDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
  `endif

    not (nD, D);

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    $width (negedge EN &&& D_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge EN, posedge D, 0, 0, notifier,,, EN_d, D_d);
    $setuphold (posedge EN, negedge D, 0, 0, notifier,,, EN_d, D_d);
  `else
    $setuphold (posedge EN, posedge D, 0, 0, notifier);
    $setuphold (posedge EN, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNQD4 (D, EN, Q);
    input D, EN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire D_d, EN_d;
        pullup (CDN);
        pullup (SDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
  `endif

    not (nD, D);

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    $width (negedge EN &&& D_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge EN, posedge D, 0, 0, notifier,,, EN_d, D_d);
    $setuphold (posedge EN, negedge D, 0, 0, notifier,,, EN_d, D_d);
  `else
    $setuphold (posedge EN, posedge D, 0, 0, notifier);
    $setuphold (posedge EN, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNSND1 (D, EN, SDN, Q, QN);
    input D, EN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, EN_d;
        pullup (CDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
  `endif

    not (nD, D);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);

  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    if (D == 1'b1 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    if (D == 1'b1 && EN == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge EN &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nD_EN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0, notifier);
      $hold (posedge EN &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0, notifier);
    $hold (posedge EN &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNSND2 (D, EN, SDN, Q, QN);
    input D, EN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, EN_d;
        pullup (CDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
  `endif

    not (nD, D);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);

  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    if (D == 1'b1 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    if (D == 1'b1 && EN == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge EN &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nD_EN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0, notifier);
      $hold (posedge EN &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0, notifier);
    $hold (posedge EN &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNSND4 (D, EN, SDN, Q, QN);
    input D, EN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, EN_d;
        pullup (CDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
  `endif

    not (nD, D);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);

  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    if (D == 1'b1 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    if (D == 1'b1 && EN == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge EN &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nD_EN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0, notifier);
      $hold (posedge EN &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0, notifier);
    $hold (posedge EN &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNSNQD1 (D, EN, SDN, Q);
    input D, EN, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, EN_d;
        pullup (CDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
  `endif

    not (nD, D);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);

  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    if (D == 1'b1 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (negedge EN &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nD_EN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0, notifier);
      $hold (posedge EN &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0, notifier);
    $hold (posedge EN &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNSNQD2 (D, EN, SDN, Q);
    input D, EN, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, EN_d;
        pullup (CDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
  `endif

    not (nD, D);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);

  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    if (D == 1'b1 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (negedge EN &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nD_EN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0, notifier);
      $hold (posedge EN &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0, notifier);
    $hold (posedge EN &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNSNQD4 (D, EN, SDN, Q);
    input D, EN, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, EN_d;
        pullup (CDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
  `endif

    not (nD, D);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);

  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    if (D == 1'b1 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (negedge EN &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nD_EN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0, notifier);
      $hold (posedge EN &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0, notifier);
    $hold (posedge EN &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module MAOI222D0 (A, B, C, ZN);
    input A, B, C;
    output ZN;
    and (I0_out, A, B);
    and (I1_out, B, C);
    and (I2_out, A, C);
    or (I3_out, I0_out, I1_out, I2_out);
    not (ZN, I3_out);

  specify
    if (B == 1'b1 && C == 1'b0)
    (A => ZN) = (0, 0);
    if (B == 1'b0 && C == 1'b1)
    (A => ZN) = (0, 0);
    if (A == 1'b1 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A == 1'b0 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MAOI222D1 (A, B, C, ZN);
    input A, B, C;
    output ZN;
    and (I0_out, A, B);
    and (I1_out, B, C);
    and (I2_out, A, C);
    or (I3_out, I0_out, I1_out, I2_out);
    not (ZN, I3_out);

  specify
    if (B == 1'b1 && C == 1'b0)
    (A => ZN) = (0, 0);
    if (B == 1'b0 && C == 1'b1)
    (A => ZN) = (0, 0);
    if (A == 1'b1 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A == 1'b0 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MAOI222D2 (A, B, C, ZN);
    input A, B, C;
    output ZN;
    and (I0_out, A, B);
    and (I1_out, B, C);
    and (I2_out, A, C);
    or (I3_out, I0_out, I1_out, I2_out);
    not (ZN, I3_out);

  specify
    if (B == 1'b1 && C == 1'b0)
    (A => ZN) = (0, 0);
    if (B == 1'b0 && C == 1'b1)
    (A => ZN) = (0, 0);
    if (A == 1'b1 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A == 1'b0 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MAOI222D4 (A, B, C, ZN);
    input A, B, C;
    output ZN;
    and (I0_out, A, B);
    and (I1_out, B, C);
    and (I2_out, A, C);
    or (I3_out, I0_out, I1_out, I2_out);
    not (ZN, I3_out);

  specify
    if (B == 1'b1 && C == 1'b0)
    (A => ZN) = (0, 0);
    if (B == 1'b0 && C == 1'b1)
    (A => ZN) = (0, 0);
    if (A == 1'b1 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A == 1'b0 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MAOI22D0 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and (I0_out, A1, A2);
    not (I1_out, I0_out);
    or (I2_out, B1, B2);
    and (ZN, I1_out, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MAOI22D1 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and (I0_out, A1, A2);
    not (I1_out, I0_out);
    or (I2_out, B1, B2);
    and (ZN, I1_out, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MAOI22D2 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and (I0_out, A1, A2);
    not (I1_out, I0_out);
    or (I2_out, B1, B2);
    and (ZN, I1_out, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MAOI22D4 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and (I0_out, A1, A2);
    not (I1_out, I0_out);
    or (I2_out, B1, B2);
    and (ZN, I1_out, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MOAI22D0 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or (I0_out, A1, A2);
    not (I1_out, I0_out);
    and (I2_out, B1, B2);
    or (ZN, I1_out, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MOAI22D1 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or (I0_out, A1, A2);
    not (I1_out, I0_out);
    and (I2_out, B1, B2);
    or (ZN, I1_out, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MOAI22D2 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or (I0_out, A1, A2);
    not (I1_out, I0_out);
    and (I2_out, B1, B2);
    or (ZN, I1_out, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MOAI22D4 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or (I0_out, A1, A2);
    not (I1_out, I0_out);
    and (I2_out, B1, B2);
    or (ZN, I1_out, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX2D0 (I0, I1, S, Z);
    input I0, I1, S;
    output Z;
    tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX2D1 (I0, I1, S, Z);
    input I0, I1, S;
    output Z;
    tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX2D2 (I0, I1, S, Z);
    input I0, I1, S;
    output Z;
    tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX2D4 (I0, I1, S, Z);
    input I0, I1, S;
    output Z;
    tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX2ND0 (I0, I1, S, ZN);
    input I0, I1, S;
    output ZN;
    tsmc_mux (I0_out, I0, I1, S);
    not (ZN, I0_out);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX2ND1 (I0, I1, S, ZN);
    input I0, I1, S;
    output ZN;
    tsmc_mux (I0_out, I0, I1, S);
    not (ZN, I0_out);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX2ND2 (I0, I1, S, ZN);
    input I0, I1, S;
    output ZN;
    tsmc_mux (I0_out, I0, I1, S);
    not (ZN, I0_out);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX2ND4 (I0, I1, S, ZN);
    input I0, I1, S;
    output ZN;
    tsmc_mux (I0_out, I0, I1, S);
    not (ZN, I0_out);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX3D0 (I0, I1, I2, S0, S1, Z);
    input I0, I1, I2, S0, S1;
    output Z;
    tsmc_mux (I0_out, I0, I1, S0);
    tsmc_mux (Z, I0_out, I2, S1);

  specify
    if (I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX3D1 (I0, I1, I2, S0, S1, Z);
    input I0, I1, I2, S0, S1;
    output Z;
    tsmc_mux (I0_out, I0, I1, S0);
    tsmc_mux (Z, I0_out, I2, S1);

  specify
    if (I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX3D2 (I0, I1, I2, S0, S1, Z);
    input I0, I1, I2, S0, S1;
    output Z;
    tsmc_mux (I0_out, I0, I1, S0);
    tsmc_mux (Z, I0_out, I2, S1);

  specify
    if (I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX3D4 (I0, I1, I2, S0, S1, Z);
    input I0, I1, I2, S0, S1;
    output Z;
    tsmc_mux (I0_out, I0, I1, S0);
    tsmc_mux (Z, I0_out, I2, S1);

  specify
    if (I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX3ND0 (I0, I1, I2, S0, S1, ZN);
    input I0, I1, I2, S0, S1;
    output ZN;
    tsmc_mux (I0_out, I0, I1, S0);
    tsmc_mux (I1_out, I0_out, I2, S1);
    not (ZN, I1_out);

  specify
    if (I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX3ND1 (I0, I1, I2, S0, S1, ZN);
    input I0, I1, I2, S0, S1;
    output ZN;
    tsmc_mux (I0_out, I0, I1, S0);
    tsmc_mux (I1_out, I0_out, I2, S1);
    not (ZN, I1_out);

  specify
    if (I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX3ND2 (I0, I1, I2, S0, S1, ZN);
    input I0, I1, I2, S0, S1;
    output ZN;
    tsmc_mux (I0_out, I0, I1, S0);
    tsmc_mux (I1_out, I0_out, I2, S1);
    not (ZN, I1_out);

  specify
    if (I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX3ND4 (I0, I1, I2, S0, S1, ZN);
    input I0, I1, I2, S0, S1;
    output ZN;
    tsmc_mux (I0_out, I0, I1, S0);
    tsmc_mux (I1_out, I0_out, I2, S1);
    not (ZN, I1_out);

  specify
    if (I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX4D0 (I0, I1, I2, I3, S0, S1, Z);
    input I0, I1, I2, I3, S0, S1;
    output Z;
    tsmc_mux (I0_out, I0, I1, S0);
    tsmc_mux (I1_out, I2, I3, S0);
    tsmc_mux (Z, I0_out, I1_out, S1);

  specify
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX4D1 (I0, I1, I2, I3, S0, S1, Z);
    input I0, I1, I2, I3, S0, S1;
    output Z;
    tsmc_mux (I0_out, I0, I1, S0);
    tsmc_mux (I1_out, I2, I3, S0);
    tsmc_mux (Z, I0_out, I1_out, S1);

  specify
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX4D2 (I0, I1, I2, I3, S0, S1, Z);
    input I0, I1, I2, I3, S0, S1;
    output Z;
    tsmc_mux (I0_out, I0, I1, S0);
    tsmc_mux (I1_out, I2, I3, S0);
    tsmc_mux (Z, I0_out, I1_out, S1);

  specify
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX4D4 (I0, I1, I2, I3, S0, S1, Z);
    input I0, I1, I2, I3, S0, S1;
    output Z;
    tsmc_mux (I0_out, I0, I1, S0);
    tsmc_mux (I1_out, I2, I3, S0);
    tsmc_mux (Z, I0_out, I1_out, S1);

  specify
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX4ND0 (I0, I1, I2, I3, S0, S1, ZN);
    input I0, I1, I2, I3, S0, S1;
    output ZN;
    tsmc_mux (I0_out, I0, I1, S0);
    tsmc_mux (I1_out, I2, I3, S0);
    tsmc_mux (I2_out, I0_out, I1_out, S1);
    not (ZN, I2_out);

  specify
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX4ND1 (I0, I1, I2, I3, S0, S1, ZN);
    input I0, I1, I2, I3, S0, S1;
    output ZN;
    tsmc_mux (I0_out, I0, I1, S0);
    tsmc_mux (I1_out, I2, I3, S0);
    tsmc_mux (I2_out, I0_out, I1_out, S1);
    not (ZN, I2_out);

  specify
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX4ND2 (I0, I1, I2, I3, S0, S1, ZN);
    input I0, I1, I2, I3, S0, S1;
    output ZN;
    tsmc_mux (I0_out, I0, I1, S0);
    tsmc_mux (I1_out, I2, I3, S0);
    tsmc_mux (I2_out, I0_out, I1_out, S1);
    not (ZN, I2_out);

  specify
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX4ND4 (I0, I1, I2, I3, S0, S1, ZN);
    input I0, I1, I2, I3, S0, S1;
    output ZN;
    tsmc_mux (I0_out, I0, I1, S0);
    tsmc_mux (I1_out, I2, I3, S0);
    tsmc_mux (I2_out, I0_out, I1_out, S1);
    not (ZN, I2_out);

  specify
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND2D0 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND2D1 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND2D2 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND2D3 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND2D4 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND2D8 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND3D0 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    and (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND3D1 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    and (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND3D2 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    and (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND3D3 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    and (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND3D4 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    and (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND3D8 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    and (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND4D0 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    and (I0_out, A1, A2, A3, A4);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND4D1 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    and (I0_out, A1, A2, A3, A4);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND4D2 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    and (I0_out, A1, A2, A3, A4);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND4D3 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    and (I0_out, A1, A2, A3, A4);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND4D4 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    and (I0_out, A1, A2, A3, A4);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND4D8 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    and (I0_out, A1, A2, A3, A4);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2D0 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    or (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2D1 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    or (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2D2 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    or (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2D3 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    or (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2D4 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    or (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2D8 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    or (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2XD0 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    or (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2XD1 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    or (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2XD2 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    or (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2XD3 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    or (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2XD4 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    or (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2XD8 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    or (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR3D0 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    or (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR3D1 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    or (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR3D2 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    or (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR3D3 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    or (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR3D4 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    or (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR3D8 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    or (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR4D0 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    or (I0_out, A1, A2, A3, A4);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR4D1 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    or (I0_out, A1, A2, A3, A4);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR4D2 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    or (I0_out, A1, A2, A3, A4);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR4D3 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    or (I0_out, A1, A2, A3, A4);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR4D4 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    or (I0_out, A1, A2, A3, A4);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR4D8 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    or (I0_out, A1, A2, A3, A4);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA211D0 (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
    or (I0_out, A1, A2);
    and (Z, I0_out, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && C == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b1)
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA211D1 (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
    or (I0_out, A1, A2);
    and (Z, I0_out, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && C == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b1)
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA211D2 (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
    or (I0_out, A1, A2);
    and (Z, I0_out, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && C == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b1)
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA211D4 (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
    or (I0_out, A1, A2);
    and (Z, I0_out, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && C == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b1)
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA21D0 (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
    or (I0_out, A1, A2);
    and (Z, I0_out, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA21D1 (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
    or (I0_out, A1, A2);
    and (Z, I0_out, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA21D2 (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
    or (I0_out, A1, A2);
    and (Z, I0_out, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA21D4 (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
    or (I0_out, A1, A2);
    and (Z, I0_out, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA221D0 (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (Z, I0_out, I1_out, C);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA221D1 (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (Z, I0_out, I1_out, C);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA221D2 (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (Z, I0_out, I1_out, C);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA221D4 (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (Z, I0_out, I1_out, C);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA222D0 (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    or (I2_out, C1, C2);
    and (Z, I0_out, I1_out, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA222D1 (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    or (I2_out, C1, C2);
    and (Z, I0_out, I1_out, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA222D2 (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    or (I2_out, C1, C2);
    and (Z, I0_out, I1_out, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA222D4 (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    or (I2_out, C1, C2);
    and (Z, I0_out, I1_out, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA22D0 (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA22D1 (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA22D2 (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA22D4 (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA31D0 (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
    or (I0_out, A1, A2, A3);
    and (Z, I0_out, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA31D1 (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
    or (I0_out, A1, A2, A3);
    and (Z, I0_out, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA31D2 (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
    or (I0_out, A1, A2, A3);
    and (Z, I0_out, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA31D4 (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
    or (I0_out, A1, A2, A3);
    and (Z, I0_out, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA32D0 (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
    or (I0_out, A1, A2, A3);
    or (I1_out, B1, B2);
    and (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA32D1 (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
    or (I0_out, A1, A2, A3);
    or (I1_out, B1, B2);
    and (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA32D2 (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
    or (I0_out, A1, A2, A3);
    or (I1_out, B1, B2);
    and (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA32D4 (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
    or (I0_out, A1, A2, A3);
    or (I1_out, B1, B2);
    and (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA33D0 (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
    or (I0_out, A1, A2, A3);
    or (I1_out, B1, B2, B3);
    and (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA33D1 (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
    or (I0_out, A1, A2, A3);
    or (I1_out, B1, B2, B3);
    and (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA33D2 (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
    or (I0_out, A1, A2, A3);
    or (I1_out, B1, B2, B3);
    and (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA33D4 (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
    or (I0_out, A1, A2, A3);
    or (I1_out, B1, B2, B3);
    and (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI211D0 (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    or (I0_out, A1, A2);
    and (I1_out, I0_out, B, C);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b1)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI211D1 (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    or (I0_out, A1, A2);
    and (I1_out, I0_out, B, C);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b1)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI211D2 (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    or (I0_out, A1, A2);
    and (I1_out, I0_out, B, C);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b1)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI211D4 (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    or (I0_out, A1, A2);
    and (I1_out, I0_out, B, C);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b1)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI21D0 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    or (I0_out, A1, A2);
    and (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI21D1 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    or (I0_out, A1, A2);
    and (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI21D2 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    or (I0_out, A1, A2);
    and (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI21D4 (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    or (I0_out, A1, A2);
    and (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI221D0 (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (I2_out, I0_out, I1_out, C);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI221D1 (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (I2_out, I0_out, I1_out, C);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI221D2 (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (I2_out, I0_out, I1_out, C);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI221D4 (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (I2_out, I0_out, I1_out, C);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI221XD4 (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (I2_out, I0_out, I1_out, C);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI222D0 (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    or (I2_out, C1, C2);
    and (I3_out, I0_out, I1_out, I2_out);
    not (ZN, I3_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI222D1 (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    or (I2_out, C1, C2);
    and (I3_out, I0_out, I1_out, I2_out);
    not (ZN, I3_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI222D2 (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    or (I2_out, C1, C2);
    and (I3_out, I0_out, I1_out, I2_out);
    not (ZN, I3_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI222D4 (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    or (I2_out, C1, C2);
    and (I3_out, I0_out, I1_out, I2_out);
    not (ZN, I3_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI222XD4 (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    or (I2_out, C1, C2);
    and (I3_out, I0_out, I1_out, I2_out);
    not (ZN, I3_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI22D0 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI22D1 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI22D2 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI22D4 (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI31D0 (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
    or (I0_out, A1, A2, A3);
    and (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI31D1 (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
    or (I0_out, A1, A2, A3);
    and (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI31D2 (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
    or (I0_out, A1, A2, A3);
    and (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI31D4 (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
    or (I0_out, A1, A2, A3);
    and (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI32D0 (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
    or (I0_out, A1, A2, A3);
    or (I1_out, B1, B2);
    and (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI32D1 (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
    or (I0_out, A1, A2, A3);
    or (I1_out, B1, B2);
    and (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI32D2 (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
    or (I0_out, A1, A2, A3);
    or (I1_out, B1, B2);
    and (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI32D4 (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
    or (I0_out, A1, A2, A3);
    or (I1_out, B1, B2);
    and (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI32XD4 (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
    or (I0_out, A1, A2, A3);
    or (I1_out, B1, B2);
    and (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI33D0 (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
    or (I0_out, A1, A2, A3);
    or (I1_out, B1, B2, B3);
    and (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI33D1 (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
    or (I0_out, A1, A2, A3);
    or (I1_out, B1, B2, B3);
    and (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI33D2 (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
    or (I0_out, A1, A2, A3);
    or (I1_out, B1, B2, B3);
    and (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI33D4 (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
    or (I0_out, A1, A2, A3);
    or (I1_out, B1, B2, B3);
    and (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI33XD4 (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
    or (I0_out, A1, A2, A3);
    or (I1_out, B1, B2, B3);
    and (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR2D0 (A1, A2, Z);
    input A1, A2;
    output Z;
    or (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR2D1 (A1, A2, Z);
    input A1, A2;
    output Z;
    or (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR2D2 (A1, A2, Z);
    input A1, A2;
    output Z;
    or (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR2D4 (A1, A2, Z);
    input A1, A2;
    output Z;
    or (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR2D8 (A1, A2, Z);
    input A1, A2;
    output Z;
    or (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR2XD1 (A1, A2, Z);
    input A1, A2;
    output Z;
    or (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR3D0 (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    or (Z, A1, A2, A3);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR3D1 (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    or (Z, A1, A2, A3);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR3D2 (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    or (Z, A1, A2, A3);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR3D4 (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    or (Z, A1, A2, A3);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR3D8 (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    or (Z, A1, A2, A3);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR3XD1 (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    or (Z, A1, A2, A3);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR4D0 (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    or (Z, A1, A2, A3, A4);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR4D1 (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    or (Z, A1, A2, A3, A4);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR4D2 (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    or (Z, A1, A2, A3, A4);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR4D4 (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    or (Z, A1, A2, A3, A4);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR4D8 (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    or (Z, A1, A2, A3, A4);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR4XD1 (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    or (Z, A1, A2, A3, A4);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module SDF4CQD0 (SI, D, SE, CP, Q);
    input SI, D, SE, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CP_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDF4CQD1 (SI, D, SE, CP, Q);
    input SI, D, SE, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CP_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDF4CQD2 (SI, D, SE, CP, Q);
    input SI, D, SE, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CP_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDF4CQD4 (SI, D, SE, CP, Q);
    input SI, D, SE, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CP_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCND0 (SI, D, SE, CP, CDN, Q, QN);
    input SI, D, SE, CP, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
  `endif
  and  (D_check, CDN_i, SE_int_not);
  buf  (CP_check, CDN_i);
  buf  (SE_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCND1 (SI, D, SE, CP, CDN, Q, QN);
    input SI, D, SE, CP, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
  `endif
  and  (D_check, CDN_i, SE_int_not);
  buf  (CP_check, CDN_i);
  buf  (SE_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCND2 (SI, D, SE, CP, CDN, Q, QN);
    input SI, D, SE, CP, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
  `endif
  and  (D_check, CDN_i, SE_int_not);
  buf  (CP_check, CDN_i);
  buf  (SE_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCND4 (SI, D, SE, CP, CDN, Q, QN);
    input SI, D, SE, CP, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
  `endif
  and  (D_check, CDN_i, SE_int_not);
  buf  (CP_check, CDN_i);
  buf  (SE_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCNQD0 (SI, D, SE, CP, CDN, Q);
    input SI, D, SE, CP, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
  `endif
  and  (D_check, CDN_i, SE_int_not);
  buf  (CP_check, CDN_i);
  buf  (SE_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCNQD1 (SI, D, SE, CP, CDN, Q);
    input SI, D, SE, CP, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
  `endif
  and  (D_check, CDN_i, SE_int_not);
  buf  (CP_check, CDN_i);
  buf  (SE_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCNQD2 (SI, D, SE, CP, CDN, Q);
    input SI, D, SE, CP, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
  `endif
  and  (D_check, CDN_i, SE_int_not);
  buf  (CP_check, CDN_i);
  buf  (SE_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCNQD4 (SI, D, SE, CP, CDN, Q);
    input SI, D, SE, CP, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
  `endif
  and  (D_check, CDN_i, SE_int_not);
  buf  (CP_check, CDN_i);
  buf  (SE_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCSND0 (SI, D, SE, CP, CDN, SDN, Q, QN);
    input SI, D, SE, CP, CDN, SDN;
    output Q, QN;
    reg notifier;
    reg flag;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SDN_SE_SI_SDFCHK, CP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_SE_nSI_SDFCHK, CP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_SI_SDFCHK, CP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_nSI_SDFCHK, CP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_SI_SDFCHK, CP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_nSI_SDFCHK, CP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_SI_SDFCHK, CP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_nSI_SDFCHK, CP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_SI_SDFCHK, nCP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_nSI_SDFCHK, nCP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_SI_SDFCHK, nCP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_nSI_SDFCHK, nCP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_SI_SDFCHK, nCP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_nSI_SDFCHK, nCP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_SI_SDFCHK, nCP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_nSI_SDFCHK, nCP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SI_SDFCHK, CDN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_SI_SDFCHK, CDN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_nSI_SDFCHK, CDN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SI_SDFCHK, CDN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_nSI_SDFCHK, CDN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_nSI_SDFCHK, CDN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_SI_SDFCHK, CDN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_nSI_SDFCHK, CDN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_SI_SDFCHK, CDN_CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_nSI_SDFCHK, CDN_CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_SI_SDFCHK, CDN_CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_nSI_SDFCHK, CDN_CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_SI_SDFCHK, CDN_CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_nSI_SDFCHK, CDN_CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_SI_SDFCHK, CDN_CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_nSI_SDFCHK, CDN_CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_SI_SDFCHK, CDN_nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_SI_SDFCHK, CDN_nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_nSI_SDFCHK, CDN_nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_SI_SDFCHK, CDN_nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_nSI_SDFCHK, CDN_nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_nSI_SDFCHK, CDN_nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_SI_SDFCHK, CDN_nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_nSI_SDFCHK, CDN_nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_SI_SDFCHK, CDN_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_nSI_SDFCHK, CDN_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SI_SDFCHK, CDN_nD_SDN_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSI_SDFCHK, CDN_D_SDN_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SDFCHK, CDN_D_SDN_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SDFCHK, CDN_nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SDN_SE_SI, CP, D, SDN, SE, SI);
    and (CP_D_SDN_SE_nSI, CP, D, SDN, SE, nSI);
    and (CP_D_SDN_nSE_SI, CP, D, SDN, nSE, SI);
    and (CP_D_SDN_nSE_nSI, CP, D, SDN, nSE, nSI);
    and (CP_nD_SDN_SE_SI, CP, nD, SDN, SE, SI);
    and (CP_nD_SDN_SE_nSI, CP, nD, SDN, SE, nSI);
    and (CP_nD_SDN_nSE_SI, CP, nD, SDN, nSE, SI);
    and (CP_nD_SDN_nSE_nSI, CP, nD, SDN, nSE, nSI);
    and (nCP_D_SDN_SE_SI, nCP, D, SDN, SE, SI);
    and (nCP_D_SDN_SE_nSI, nCP, D, SDN, SE, nSI);
    and (nCP_D_SDN_nSE_SI, nCP, D, SDN, nSE, SI);
    and (nCP_D_SDN_nSE_nSI, nCP, D, SDN, nSE, nSI);
    and (nCP_nD_SDN_SE_SI, nCP, nD, SDN, SE, SI);
    and (nCP_nD_SDN_SE_nSI, nCP, nD, SDN, SE, nSI);
    and (nCP_nD_SDN_nSE_SI, nCP, nD, SDN, nSE, SI);
    and (nCP_nD_SDN_nSE_nSI, nCP, nD, SDN, nSE, nSI);
    and (CDN_D_SDN_SE_SI, CDN, D, SDN, SE, SI);
    and (CDN_D_SDN_nSE_SI, CDN, D, SDN, nSE, SI);
    and (CDN_D_SDN_nSE_nSI, CDN, D, SDN, nSE, nSI);
    and (CDN_nD_SDN_SE_SI, CDN, nD, SDN, SE, SI);
    and (CDN_D_SDN_SE_nSI, CDN, D, SDN, SE, nSI);
    and (CDN_nD_SDN_SE_nSI, CDN, nD, SDN, SE, nSI);
    and (CDN_nD_SDN_nSE_SI, CDN, nD, SDN, nSE, SI);
    and (CDN_nD_SDN_nSE_nSI, CDN, nD, SDN, nSE, nSI);
    and (CDN_CP_D_SE_SI, CDN, CP, D, SE, SI);
    and (CDN_CP_D_SE_nSI, CDN, CP, D, SE, nSI);
    and (CDN_CP_D_nSE_SI, CDN, CP, D, nSE, SI);
    and (CDN_CP_D_nSE_nSI, CDN, CP, D, nSE, nSI);
    and (CDN_CP_nD_SE_SI, CDN, CP, nD, SE, SI);
    and (CDN_CP_nD_SE_nSI, CDN, CP, nD, SE, nSI);
    and (CDN_CP_nD_nSE_SI, CDN, CP, nD, nSE, SI);
    and (CDN_CP_nD_nSE_nSI, CDN, CP, nD, nSE, nSI);
    and (CDN_nCP_D_SE_SI, CDN, nCP, D, SE, SI);
    and (CDN_nCP_D_nSE_SI, CDN, nCP, D, nSE, SI);
    and (CDN_nCP_D_nSE_nSI, CDN, nCP, D, nSE, nSI);
    and (CDN_nCP_nD_SE_SI, CDN, nCP, nD, SE, SI);
    and (CDN_nCP_D_SE_nSI, CDN, nCP, D, SE, nSI);
    and (CDN_nCP_nD_SE_nSI, CDN, nCP, nD, SE, nSI);
    and (CDN_nCP_nD_nSE_SI, CDN, nCP, nD, nSE, SI);
    and (CDN_nCP_nD_nSE_nSI, CDN, nCP, nD, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_SDN_nSE_SI, CDN, SDN, nSE, SI);
    and (CDN_SDN_nSE_nSI, CDN, SDN, nSE, nSI);
    and (CDN_nD_SDN_SI, CDN, nD, SDN, SI);
    and (CDN_D_SDN_nSI, CDN, D, SDN, nSI);
    and (CDN_D_SDN_SE, CDN, D, SDN, SE);
    and (CDN_nD_SDN_SE, CDN, nD, SDN, SE);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SDN_i, SE);
  `endif
  and  (D_check, CDN_i, SDN_i, SE_int_not);
  and  (CP_check, CDN_i, SDN_i);
  and  (SE_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCSND1 (SI, D, SE, CP, CDN, SDN, Q, QN);
    input SI, D, SE, CP, CDN, SDN;
    output Q, QN;
    reg notifier;
    reg flag;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SDN_SE_SI_SDFCHK, CP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_SE_nSI_SDFCHK, CP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_SI_SDFCHK, CP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_nSI_SDFCHK, CP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_SI_SDFCHK, CP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_nSI_SDFCHK, CP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_SI_SDFCHK, CP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_nSI_SDFCHK, CP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_SI_SDFCHK, nCP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_nSI_SDFCHK, nCP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_SI_SDFCHK, nCP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_nSI_SDFCHK, nCP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_SI_SDFCHK, nCP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_nSI_SDFCHK, nCP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_SI_SDFCHK, nCP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_nSI_SDFCHK, nCP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SI_SDFCHK, CDN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_SI_SDFCHK, CDN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_nSI_SDFCHK, CDN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SI_SDFCHK, CDN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_nSI_SDFCHK, CDN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_nSI_SDFCHK, CDN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_SI_SDFCHK, CDN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_nSI_SDFCHK, CDN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_SI_SDFCHK, CDN_CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_nSI_SDFCHK, CDN_CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_SI_SDFCHK, CDN_CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_nSI_SDFCHK, CDN_CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_SI_SDFCHK, CDN_CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_nSI_SDFCHK, CDN_CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_SI_SDFCHK, CDN_CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_nSI_SDFCHK, CDN_CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_SI_SDFCHK, CDN_nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_SI_SDFCHK, CDN_nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_nSI_SDFCHK, CDN_nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_SI_SDFCHK, CDN_nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_nSI_SDFCHK, CDN_nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_nSI_SDFCHK, CDN_nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_SI_SDFCHK, CDN_nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_nSI_SDFCHK, CDN_nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_SI_SDFCHK, CDN_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_nSI_SDFCHK, CDN_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SI_SDFCHK, CDN_nD_SDN_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSI_SDFCHK, CDN_D_SDN_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SDFCHK, CDN_D_SDN_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SDFCHK, CDN_nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SDN_SE_SI, CP, D, SDN, SE, SI);
    and (CP_D_SDN_SE_nSI, CP, D, SDN, SE, nSI);
    and (CP_D_SDN_nSE_SI, CP, D, SDN, nSE, SI);
    and (CP_D_SDN_nSE_nSI, CP, D, SDN, nSE, nSI);
    and (CP_nD_SDN_SE_SI, CP, nD, SDN, SE, SI);
    and (CP_nD_SDN_SE_nSI, CP, nD, SDN, SE, nSI);
    and (CP_nD_SDN_nSE_SI, CP, nD, SDN, nSE, SI);
    and (CP_nD_SDN_nSE_nSI, CP, nD, SDN, nSE, nSI);
    and (nCP_D_SDN_SE_SI, nCP, D, SDN, SE, SI);
    and (nCP_D_SDN_SE_nSI, nCP, D, SDN, SE, nSI);
    and (nCP_D_SDN_nSE_SI, nCP, D, SDN, nSE, SI);
    and (nCP_D_SDN_nSE_nSI, nCP, D, SDN, nSE, nSI);
    and (nCP_nD_SDN_SE_SI, nCP, nD, SDN, SE, SI);
    and (nCP_nD_SDN_SE_nSI, nCP, nD, SDN, SE, nSI);
    and (nCP_nD_SDN_nSE_SI, nCP, nD, SDN, nSE, SI);
    and (nCP_nD_SDN_nSE_nSI, nCP, nD, SDN, nSE, nSI);
    and (CDN_D_SDN_SE_SI, CDN, D, SDN, SE, SI);
    and (CDN_D_SDN_nSE_SI, CDN, D, SDN, nSE, SI);
    and (CDN_D_SDN_nSE_nSI, CDN, D, SDN, nSE, nSI);
    and (CDN_nD_SDN_SE_SI, CDN, nD, SDN, SE, SI);
    and (CDN_D_SDN_SE_nSI, CDN, D, SDN, SE, nSI);
    and (CDN_nD_SDN_SE_nSI, CDN, nD, SDN, SE, nSI);
    and (CDN_nD_SDN_nSE_SI, CDN, nD, SDN, nSE, SI);
    and (CDN_nD_SDN_nSE_nSI, CDN, nD, SDN, nSE, nSI);
    and (CDN_CP_D_SE_SI, CDN, CP, D, SE, SI);
    and (CDN_CP_D_SE_nSI, CDN, CP, D, SE, nSI);
    and (CDN_CP_D_nSE_SI, CDN, CP, D, nSE, SI);
    and (CDN_CP_D_nSE_nSI, CDN, CP, D, nSE, nSI);
    and (CDN_CP_nD_SE_SI, CDN, CP, nD, SE, SI);
    and (CDN_CP_nD_SE_nSI, CDN, CP, nD, SE, nSI);
    and (CDN_CP_nD_nSE_SI, CDN, CP, nD, nSE, SI);
    and (CDN_CP_nD_nSE_nSI, CDN, CP, nD, nSE, nSI);
    and (CDN_nCP_D_SE_SI, CDN, nCP, D, SE, SI);
    and (CDN_nCP_D_nSE_SI, CDN, nCP, D, nSE, SI);
    and (CDN_nCP_D_nSE_nSI, CDN, nCP, D, nSE, nSI);
    and (CDN_nCP_nD_SE_SI, CDN, nCP, nD, SE, SI);
    and (CDN_nCP_D_SE_nSI, CDN, nCP, D, SE, nSI);
    and (CDN_nCP_nD_SE_nSI, CDN, nCP, nD, SE, nSI);
    and (CDN_nCP_nD_nSE_SI, CDN, nCP, nD, nSE, SI);
    and (CDN_nCP_nD_nSE_nSI, CDN, nCP, nD, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_SDN_nSE_SI, CDN, SDN, nSE, SI);
    and (CDN_SDN_nSE_nSI, CDN, SDN, nSE, nSI);
    and (CDN_nD_SDN_SI, CDN, nD, SDN, SI);
    and (CDN_D_SDN_nSI, CDN, D, SDN, nSI);
    and (CDN_D_SDN_SE, CDN, D, SDN, SE);
    and (CDN_nD_SDN_SE, CDN, nD, SDN, SE);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SDN_i, SE);
  `endif
  and  (D_check, CDN_i, SDN_i, SE_int_not);
  and  (CP_check, CDN_i, SDN_i);
  and  (SE_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCSND2 (SI, D, SE, CP, CDN, SDN, Q, QN);
    input SI, D, SE, CP, CDN, SDN;
    output Q, QN;
    reg notifier;
    reg flag;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SDN_SE_SI_SDFCHK, CP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_SE_nSI_SDFCHK, CP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_SI_SDFCHK, CP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_nSI_SDFCHK, CP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_SI_SDFCHK, CP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_nSI_SDFCHK, CP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_SI_SDFCHK, CP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_nSI_SDFCHK, CP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_SI_SDFCHK, nCP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_nSI_SDFCHK, nCP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_SI_SDFCHK, nCP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_nSI_SDFCHK, nCP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_SI_SDFCHK, nCP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_nSI_SDFCHK, nCP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_SI_SDFCHK, nCP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_nSI_SDFCHK, nCP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SI_SDFCHK, CDN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_SI_SDFCHK, CDN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_nSI_SDFCHK, CDN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SI_SDFCHK, CDN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_nSI_SDFCHK, CDN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_nSI_SDFCHK, CDN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_SI_SDFCHK, CDN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_nSI_SDFCHK, CDN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_SI_SDFCHK, CDN_CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_nSI_SDFCHK, CDN_CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_SI_SDFCHK, CDN_CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_nSI_SDFCHK, CDN_CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_SI_SDFCHK, CDN_CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_nSI_SDFCHK, CDN_CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_SI_SDFCHK, CDN_CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_nSI_SDFCHK, CDN_CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_SI_SDFCHK, CDN_nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_SI_SDFCHK, CDN_nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_nSI_SDFCHK, CDN_nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_SI_SDFCHK, CDN_nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_nSI_SDFCHK, CDN_nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_nSI_SDFCHK, CDN_nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_SI_SDFCHK, CDN_nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_nSI_SDFCHK, CDN_nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_SI_SDFCHK, CDN_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_nSI_SDFCHK, CDN_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SI_SDFCHK, CDN_nD_SDN_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSI_SDFCHK, CDN_D_SDN_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SDFCHK, CDN_D_SDN_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SDFCHK, CDN_nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SDN_SE_SI, CP, D, SDN, SE, SI);
    and (CP_D_SDN_SE_nSI, CP, D, SDN, SE, nSI);
    and (CP_D_SDN_nSE_SI, CP, D, SDN, nSE, SI);
    and (CP_D_SDN_nSE_nSI, CP, D, SDN, nSE, nSI);
    and (CP_nD_SDN_SE_SI, CP, nD, SDN, SE, SI);
    and (CP_nD_SDN_SE_nSI, CP, nD, SDN, SE, nSI);
    and (CP_nD_SDN_nSE_SI, CP, nD, SDN, nSE, SI);
    and (CP_nD_SDN_nSE_nSI, CP, nD, SDN, nSE, nSI);
    and (nCP_D_SDN_SE_SI, nCP, D, SDN, SE, SI);
    and (nCP_D_SDN_SE_nSI, nCP, D, SDN, SE, nSI);
    and (nCP_D_SDN_nSE_SI, nCP, D, SDN, nSE, SI);
    and (nCP_D_SDN_nSE_nSI, nCP, D, SDN, nSE, nSI);
    and (nCP_nD_SDN_SE_SI, nCP, nD, SDN, SE, SI);
    and (nCP_nD_SDN_SE_nSI, nCP, nD, SDN, SE, nSI);
    and (nCP_nD_SDN_nSE_SI, nCP, nD, SDN, nSE, SI);
    and (nCP_nD_SDN_nSE_nSI, nCP, nD, SDN, nSE, nSI);
    and (CDN_D_SDN_SE_SI, CDN, D, SDN, SE, SI);
    and (CDN_D_SDN_nSE_SI, CDN, D, SDN, nSE, SI);
    and (CDN_D_SDN_nSE_nSI, CDN, D, SDN, nSE, nSI);
    and (CDN_nD_SDN_SE_SI, CDN, nD, SDN, SE, SI);
    and (CDN_D_SDN_SE_nSI, CDN, D, SDN, SE, nSI);
    and (CDN_nD_SDN_SE_nSI, CDN, nD, SDN, SE, nSI);
    and (CDN_nD_SDN_nSE_SI, CDN, nD, SDN, nSE, SI);
    and (CDN_nD_SDN_nSE_nSI, CDN, nD, SDN, nSE, nSI);
    and (CDN_CP_D_SE_SI, CDN, CP, D, SE, SI);
    and (CDN_CP_D_SE_nSI, CDN, CP, D, SE, nSI);
    and (CDN_CP_D_nSE_SI, CDN, CP, D, nSE, SI);
    and (CDN_CP_D_nSE_nSI, CDN, CP, D, nSE, nSI);
    and (CDN_CP_nD_SE_SI, CDN, CP, nD, SE, SI);
    and (CDN_CP_nD_SE_nSI, CDN, CP, nD, SE, nSI);
    and (CDN_CP_nD_nSE_SI, CDN, CP, nD, nSE, SI);
    and (CDN_CP_nD_nSE_nSI, CDN, CP, nD, nSE, nSI);
    and (CDN_nCP_D_SE_SI, CDN, nCP, D, SE, SI);
    and (CDN_nCP_D_nSE_SI, CDN, nCP, D, nSE, SI);
    and (CDN_nCP_D_nSE_nSI, CDN, nCP, D, nSE, nSI);
    and (CDN_nCP_nD_SE_SI, CDN, nCP, nD, SE, SI);
    and (CDN_nCP_D_SE_nSI, CDN, nCP, D, SE, nSI);
    and (CDN_nCP_nD_SE_nSI, CDN, nCP, nD, SE, nSI);
    and (CDN_nCP_nD_nSE_SI, CDN, nCP, nD, nSE, SI);
    and (CDN_nCP_nD_nSE_nSI, CDN, nCP, nD, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_SDN_nSE_SI, CDN, SDN, nSE, SI);
    and (CDN_SDN_nSE_nSI, CDN, SDN, nSE, nSI);
    and (CDN_nD_SDN_SI, CDN, nD, SDN, SI);
    and (CDN_D_SDN_nSI, CDN, D, SDN, nSI);
    and (CDN_D_SDN_SE, CDN, D, SDN, SE);
    and (CDN_nD_SDN_SE, CDN, nD, SDN, SE);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SDN_i, SE);
  `endif
  and  (D_check, CDN_i, SDN_i, SE_int_not);
  and  (CP_check, CDN_i, SDN_i);
  and  (SE_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCSND4 (SI, D, SE, CP, CDN, SDN, Q, QN);
    input SI, D, SE, CP, CDN, SDN;
    output Q, QN;
    reg notifier;
    reg flag;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SDN_SE_SI_SDFCHK, CP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_SE_nSI_SDFCHK, CP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_SI_SDFCHK, CP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_nSI_SDFCHK, CP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_SI_SDFCHK, CP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_nSI_SDFCHK, CP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_SI_SDFCHK, CP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_nSI_SDFCHK, CP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_SI_SDFCHK, nCP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_nSI_SDFCHK, nCP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_SI_SDFCHK, nCP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_nSI_SDFCHK, nCP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_SI_SDFCHK, nCP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_nSI_SDFCHK, nCP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_SI_SDFCHK, nCP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_nSI_SDFCHK, nCP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SI_SDFCHK, CDN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_SI_SDFCHK, CDN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_nSI_SDFCHK, CDN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SI_SDFCHK, CDN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_nSI_SDFCHK, CDN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_nSI_SDFCHK, CDN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_SI_SDFCHK, CDN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_nSI_SDFCHK, CDN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_SI_SDFCHK, CDN_CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_nSI_SDFCHK, CDN_CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_SI_SDFCHK, CDN_CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_nSI_SDFCHK, CDN_CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_SI_SDFCHK, CDN_CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_nSI_SDFCHK, CDN_CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_SI_SDFCHK, CDN_CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_nSI_SDFCHK, CDN_CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_SI_SDFCHK, CDN_nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_SI_SDFCHK, CDN_nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_nSI_SDFCHK, CDN_nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_SI_SDFCHK, CDN_nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_nSI_SDFCHK, CDN_nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_nSI_SDFCHK, CDN_nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_SI_SDFCHK, CDN_nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_nSI_SDFCHK, CDN_nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_SI_SDFCHK, CDN_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_nSI_SDFCHK, CDN_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SI_SDFCHK, CDN_nD_SDN_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSI_SDFCHK, CDN_D_SDN_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SDFCHK, CDN_D_SDN_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SDFCHK, CDN_nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SDN_SE_SI, CP, D, SDN, SE, SI);
    and (CP_D_SDN_SE_nSI, CP, D, SDN, SE, nSI);
    and (CP_D_SDN_nSE_SI, CP, D, SDN, nSE, SI);
    and (CP_D_SDN_nSE_nSI, CP, D, SDN, nSE, nSI);
    and (CP_nD_SDN_SE_SI, CP, nD, SDN, SE, SI);
    and (CP_nD_SDN_SE_nSI, CP, nD, SDN, SE, nSI);
    and (CP_nD_SDN_nSE_SI, CP, nD, SDN, nSE, SI);
    and (CP_nD_SDN_nSE_nSI, CP, nD, SDN, nSE, nSI);
    and (nCP_D_SDN_SE_SI, nCP, D, SDN, SE, SI);
    and (nCP_D_SDN_SE_nSI, nCP, D, SDN, SE, nSI);
    and (nCP_D_SDN_nSE_SI, nCP, D, SDN, nSE, SI);
    and (nCP_D_SDN_nSE_nSI, nCP, D, SDN, nSE, nSI);
    and (nCP_nD_SDN_SE_SI, nCP, nD, SDN, SE, SI);
    and (nCP_nD_SDN_SE_nSI, nCP, nD, SDN, SE, nSI);
    and (nCP_nD_SDN_nSE_SI, nCP, nD, SDN, nSE, SI);
    and (nCP_nD_SDN_nSE_nSI, nCP, nD, SDN, nSE, nSI);
    and (CDN_D_SDN_SE_SI, CDN, D, SDN, SE, SI);
    and (CDN_D_SDN_nSE_SI, CDN, D, SDN, nSE, SI);
    and (CDN_D_SDN_nSE_nSI, CDN, D, SDN, nSE, nSI);
    and (CDN_nD_SDN_SE_SI, CDN, nD, SDN, SE, SI);
    and (CDN_D_SDN_SE_nSI, CDN, D, SDN, SE, nSI);
    and (CDN_nD_SDN_SE_nSI, CDN, nD, SDN, SE, nSI);
    and (CDN_nD_SDN_nSE_SI, CDN, nD, SDN, nSE, SI);
    and (CDN_nD_SDN_nSE_nSI, CDN, nD, SDN, nSE, nSI);
    and (CDN_CP_D_SE_SI, CDN, CP, D, SE, SI);
    and (CDN_CP_D_SE_nSI, CDN, CP, D, SE, nSI);
    and (CDN_CP_D_nSE_SI, CDN, CP, D, nSE, SI);
    and (CDN_CP_D_nSE_nSI, CDN, CP, D, nSE, nSI);
    and (CDN_CP_nD_SE_SI, CDN, CP, nD, SE, SI);
    and (CDN_CP_nD_SE_nSI, CDN, CP, nD, SE, nSI);
    and (CDN_CP_nD_nSE_SI, CDN, CP, nD, nSE, SI);
    and (CDN_CP_nD_nSE_nSI, CDN, CP, nD, nSE, nSI);
    and (CDN_nCP_D_SE_SI, CDN, nCP, D, SE, SI);
    and (CDN_nCP_D_nSE_SI, CDN, nCP, D, nSE, SI);
    and (CDN_nCP_D_nSE_nSI, CDN, nCP, D, nSE, nSI);
    and (CDN_nCP_nD_SE_SI, CDN, nCP, nD, SE, SI);
    and (CDN_nCP_D_SE_nSI, CDN, nCP, D, SE, nSI);
    and (CDN_nCP_nD_SE_nSI, CDN, nCP, nD, SE, nSI);
    and (CDN_nCP_nD_nSE_SI, CDN, nCP, nD, nSE, SI);
    and (CDN_nCP_nD_nSE_nSI, CDN, nCP, nD, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_SDN_nSE_SI, CDN, SDN, nSE, SI);
    and (CDN_SDN_nSE_nSI, CDN, SDN, nSE, nSI);
    and (CDN_nD_SDN_SI, CDN, nD, SDN, SI);
    and (CDN_D_SDN_nSI, CDN, D, SDN, nSI);
    and (CDN_D_SDN_SE, CDN, D, SDN, SE);
    and (CDN_nD_SDN_SE, CDN, nD, SDN, SE);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SDN_i, SE);
  `endif
  and  (D_check, CDN_i, SDN_i, SE_int_not);
  and  (CP_check, CDN_i, SDN_i);
  and  (SE_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCSNQD0 (SI, D, SE, CP, CDN, SDN, Q);
    input SI, D, SE, CP, CDN, SDN;
    output Q;
    reg notifier;
    reg flag;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SDN_SE_SI_SDFCHK, CP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_SE_nSI_SDFCHK, CP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_SI_SDFCHK, CP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_nSI_SDFCHK, CP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_SI_SDFCHK, CP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_nSI_SDFCHK, CP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_SI_SDFCHK, CP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_nSI_SDFCHK, CP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_SI_SDFCHK, nCP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_nSI_SDFCHK, nCP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_SI_SDFCHK, nCP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_nSI_SDFCHK, nCP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_SI_SDFCHK, nCP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_nSI_SDFCHK, nCP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_SI_SDFCHK, nCP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_nSI_SDFCHK, nCP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SI_SDFCHK, CDN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_SI_SDFCHK, CDN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_nSI_SDFCHK, CDN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SI_SDFCHK, CDN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_nSI_SDFCHK, CDN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_nSI_SDFCHK, CDN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_SI_SDFCHK, CDN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_nSI_SDFCHK, CDN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_SI_SDFCHK, CDN_CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_nSI_SDFCHK, CDN_CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_SI_SDFCHK, CDN_CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_nSI_SDFCHK, CDN_CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_SI_SDFCHK, CDN_CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_nSI_SDFCHK, CDN_CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_SI_SDFCHK, CDN_CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_nSI_SDFCHK, CDN_CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_SI_SDFCHK, CDN_nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_SI_SDFCHK, CDN_nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_nSI_SDFCHK, CDN_nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_SI_SDFCHK, CDN_nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_nSI_SDFCHK, CDN_nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_nSI_SDFCHK, CDN_nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_SI_SDFCHK, CDN_nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_nSI_SDFCHK, CDN_nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_SI_SDFCHK, CDN_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_nSI_SDFCHK, CDN_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SI_SDFCHK, CDN_nD_SDN_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSI_SDFCHK, CDN_D_SDN_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SDFCHK, CDN_D_SDN_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SDFCHK, CDN_nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SDN_SE_SI, CP, D, SDN, SE, SI);
    and (CP_D_SDN_SE_nSI, CP, D, SDN, SE, nSI);
    and (CP_D_SDN_nSE_SI, CP, D, SDN, nSE, SI);
    and (CP_D_SDN_nSE_nSI, CP, D, SDN, nSE, nSI);
    and (CP_nD_SDN_SE_SI, CP, nD, SDN, SE, SI);
    and (CP_nD_SDN_SE_nSI, CP, nD, SDN, SE, nSI);
    and (CP_nD_SDN_nSE_SI, CP, nD, SDN, nSE, SI);
    and (CP_nD_SDN_nSE_nSI, CP, nD, SDN, nSE, nSI);
    and (nCP_D_SDN_SE_SI, nCP, D, SDN, SE, SI);
    and (nCP_D_SDN_SE_nSI, nCP, D, SDN, SE, nSI);
    and (nCP_D_SDN_nSE_SI, nCP, D, SDN, nSE, SI);
    and (nCP_D_SDN_nSE_nSI, nCP, D, SDN, nSE, nSI);
    and (nCP_nD_SDN_SE_SI, nCP, nD, SDN, SE, SI);
    and (nCP_nD_SDN_SE_nSI, nCP, nD, SDN, SE, nSI);
    and (nCP_nD_SDN_nSE_SI, nCP, nD, SDN, nSE, SI);
    and (nCP_nD_SDN_nSE_nSI, nCP, nD, SDN, nSE, nSI);
    and (CDN_D_SDN_SE_SI, CDN, D, SDN, SE, SI);
    and (CDN_D_SDN_nSE_SI, CDN, D, SDN, nSE, SI);
    and (CDN_D_SDN_nSE_nSI, CDN, D, SDN, nSE, nSI);
    and (CDN_nD_SDN_SE_SI, CDN, nD, SDN, SE, SI);
    and (CDN_D_SDN_SE_nSI, CDN, D, SDN, SE, nSI);
    and (CDN_nD_SDN_SE_nSI, CDN, nD, SDN, SE, nSI);
    and (CDN_nD_SDN_nSE_SI, CDN, nD, SDN, nSE, SI);
    and (CDN_nD_SDN_nSE_nSI, CDN, nD, SDN, nSE, nSI);
    and (CDN_CP_D_SE_SI, CDN, CP, D, SE, SI);
    and (CDN_CP_D_SE_nSI, CDN, CP, D, SE, nSI);
    and (CDN_CP_D_nSE_SI, CDN, CP, D, nSE, SI);
    and (CDN_CP_D_nSE_nSI, CDN, CP, D, nSE, nSI);
    and (CDN_CP_nD_SE_SI, CDN, CP, nD, SE, SI);
    and (CDN_CP_nD_SE_nSI, CDN, CP, nD, SE, nSI);
    and (CDN_CP_nD_nSE_SI, CDN, CP, nD, nSE, SI);
    and (CDN_CP_nD_nSE_nSI, CDN, CP, nD, nSE, nSI);
    and (CDN_nCP_D_SE_SI, CDN, nCP, D, SE, SI);
    and (CDN_nCP_D_nSE_SI, CDN, nCP, D, nSE, SI);
    and (CDN_nCP_D_nSE_nSI, CDN, nCP, D, nSE, nSI);
    and (CDN_nCP_nD_SE_SI, CDN, nCP, nD, SE, SI);
    and (CDN_nCP_D_SE_nSI, CDN, nCP, D, SE, nSI);
    and (CDN_nCP_nD_SE_nSI, CDN, nCP, nD, SE, nSI);
    and (CDN_nCP_nD_nSE_SI, CDN, nCP, nD, nSE, SI);
    and (CDN_nCP_nD_nSE_nSI, CDN, nCP, nD, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_SDN_nSE_SI, CDN, SDN, nSE, SI);
    and (CDN_SDN_nSE_nSI, CDN, SDN, nSE, nSI);
    and (CDN_nD_SDN_SI, CDN, nD, SDN, SI);
    and (CDN_D_SDN_nSI, CDN, D, SDN, nSI);
    and (CDN_D_SDN_SE, CDN, D, SDN, SE);
    and (CDN_nD_SDN_SE, CDN, nD, SDN, SE);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SDN_i, SE);
  `endif
  and  (D_check, CDN_i, SDN_i, SE_int_not);
  and  (CP_check, CDN_i, SDN_i);
  and  (SE_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCSNQD1 (SI, D, SE, CP, CDN, SDN, Q);
    input SI, D, SE, CP, CDN, SDN;
    output Q;
    reg notifier;
    reg flag;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SDN_SE_SI_SDFCHK, CP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_SE_nSI_SDFCHK, CP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_SI_SDFCHK, CP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_nSI_SDFCHK, CP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_SI_SDFCHK, CP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_nSI_SDFCHK, CP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_SI_SDFCHK, CP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_nSI_SDFCHK, CP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_SI_SDFCHK, nCP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_nSI_SDFCHK, nCP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_SI_SDFCHK, nCP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_nSI_SDFCHK, nCP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_SI_SDFCHK, nCP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_nSI_SDFCHK, nCP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_SI_SDFCHK, nCP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_nSI_SDFCHK, nCP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SI_SDFCHK, CDN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_SI_SDFCHK, CDN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_nSI_SDFCHK, CDN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SI_SDFCHK, CDN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_nSI_SDFCHK, CDN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_nSI_SDFCHK, CDN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_SI_SDFCHK, CDN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_nSI_SDFCHK, CDN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_SI_SDFCHK, CDN_CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_nSI_SDFCHK, CDN_CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_SI_SDFCHK, CDN_CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_nSI_SDFCHK, CDN_CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_SI_SDFCHK, CDN_CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_nSI_SDFCHK, CDN_CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_SI_SDFCHK, CDN_CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_nSI_SDFCHK, CDN_CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_SI_SDFCHK, CDN_nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_SI_SDFCHK, CDN_nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_nSI_SDFCHK, CDN_nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_SI_SDFCHK, CDN_nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_nSI_SDFCHK, CDN_nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_nSI_SDFCHK, CDN_nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_SI_SDFCHK, CDN_nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_nSI_SDFCHK, CDN_nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_SI_SDFCHK, CDN_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_nSI_SDFCHK, CDN_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SI_SDFCHK, CDN_nD_SDN_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSI_SDFCHK, CDN_D_SDN_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SDFCHK, CDN_D_SDN_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SDFCHK, CDN_nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SDN_SE_SI, CP, D, SDN, SE, SI);
    and (CP_D_SDN_SE_nSI, CP, D, SDN, SE, nSI);
    and (CP_D_SDN_nSE_SI, CP, D, SDN, nSE, SI);
    and (CP_D_SDN_nSE_nSI, CP, D, SDN, nSE, nSI);
    and (CP_nD_SDN_SE_SI, CP, nD, SDN, SE, SI);
    and (CP_nD_SDN_SE_nSI, CP, nD, SDN, SE, nSI);
    and (CP_nD_SDN_nSE_SI, CP, nD, SDN, nSE, SI);
    and (CP_nD_SDN_nSE_nSI, CP, nD, SDN, nSE, nSI);
    and (nCP_D_SDN_SE_SI, nCP, D, SDN, SE, SI);
    and (nCP_D_SDN_SE_nSI, nCP, D, SDN, SE, nSI);
    and (nCP_D_SDN_nSE_SI, nCP, D, SDN, nSE, SI);
    and (nCP_D_SDN_nSE_nSI, nCP, D, SDN, nSE, nSI);
    and (nCP_nD_SDN_SE_SI, nCP, nD, SDN, SE, SI);
    and (nCP_nD_SDN_SE_nSI, nCP, nD, SDN, SE, nSI);
    and (nCP_nD_SDN_nSE_SI, nCP, nD, SDN, nSE, SI);
    and (nCP_nD_SDN_nSE_nSI, nCP, nD, SDN, nSE, nSI);
    and (CDN_D_SDN_SE_SI, CDN, D, SDN, SE, SI);
    and (CDN_D_SDN_nSE_SI, CDN, D, SDN, nSE, SI);
    and (CDN_D_SDN_nSE_nSI, CDN, D, SDN, nSE, nSI);
    and (CDN_nD_SDN_SE_SI, CDN, nD, SDN, SE, SI);
    and (CDN_D_SDN_SE_nSI, CDN, D, SDN, SE, nSI);
    and (CDN_nD_SDN_SE_nSI, CDN, nD, SDN, SE, nSI);
    and (CDN_nD_SDN_nSE_SI, CDN, nD, SDN, nSE, SI);
    and (CDN_nD_SDN_nSE_nSI, CDN, nD, SDN, nSE, nSI);
    and (CDN_CP_D_SE_SI, CDN, CP, D, SE, SI);
    and (CDN_CP_D_SE_nSI, CDN, CP, D, SE, nSI);
    and (CDN_CP_D_nSE_SI, CDN, CP, D, nSE, SI);
    and (CDN_CP_D_nSE_nSI, CDN, CP, D, nSE, nSI);
    and (CDN_CP_nD_SE_SI, CDN, CP, nD, SE, SI);
    and (CDN_CP_nD_SE_nSI, CDN, CP, nD, SE, nSI);
    and (CDN_CP_nD_nSE_SI, CDN, CP, nD, nSE, SI);
    and (CDN_CP_nD_nSE_nSI, CDN, CP, nD, nSE, nSI);
    and (CDN_nCP_D_SE_SI, CDN, nCP, D, SE, SI);
    and (CDN_nCP_D_nSE_SI, CDN, nCP, D, nSE, SI);
    and (CDN_nCP_D_nSE_nSI, CDN, nCP, D, nSE, nSI);
    and (CDN_nCP_nD_SE_SI, CDN, nCP, nD, SE, SI);
    and (CDN_nCP_D_SE_nSI, CDN, nCP, D, SE, nSI);
    and (CDN_nCP_nD_SE_nSI, CDN, nCP, nD, SE, nSI);
    and (CDN_nCP_nD_nSE_SI, CDN, nCP, nD, nSE, SI);
    and (CDN_nCP_nD_nSE_nSI, CDN, nCP, nD, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_SDN_nSE_SI, CDN, SDN, nSE, SI);
    and (CDN_SDN_nSE_nSI, CDN, SDN, nSE, nSI);
    and (CDN_nD_SDN_SI, CDN, nD, SDN, SI);
    and (CDN_D_SDN_nSI, CDN, D, SDN, nSI);
    and (CDN_D_SDN_SE, CDN, D, SDN, SE);
    and (CDN_nD_SDN_SE, CDN, nD, SDN, SE);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SDN_i, SE);
  `endif
  and  (D_check, CDN_i, SDN_i, SE_int_not);
  and  (CP_check, CDN_i, SDN_i);
  and  (SE_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCSNQD2 (SI, D, SE, CP, CDN, SDN, Q);
    input SI, D, SE, CP, CDN, SDN;
    output Q;
    reg notifier;
    reg flag;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SDN_SE_SI_SDFCHK, CP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_SE_nSI_SDFCHK, CP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_SI_SDFCHK, CP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_nSI_SDFCHK, CP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_SI_SDFCHK, CP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_nSI_SDFCHK, CP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_SI_SDFCHK, CP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_nSI_SDFCHK, CP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_SI_SDFCHK, nCP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_nSI_SDFCHK, nCP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_SI_SDFCHK, nCP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_nSI_SDFCHK, nCP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_SI_SDFCHK, nCP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_nSI_SDFCHK, nCP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_SI_SDFCHK, nCP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_nSI_SDFCHK, nCP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SI_SDFCHK, CDN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_SI_SDFCHK, CDN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_nSI_SDFCHK, CDN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SI_SDFCHK, CDN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_nSI_SDFCHK, CDN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_nSI_SDFCHK, CDN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_SI_SDFCHK, CDN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_nSI_SDFCHK, CDN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_SI_SDFCHK, CDN_CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_nSI_SDFCHK, CDN_CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_SI_SDFCHK, CDN_CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_nSI_SDFCHK, CDN_CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_SI_SDFCHK, CDN_CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_nSI_SDFCHK, CDN_CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_SI_SDFCHK, CDN_CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_nSI_SDFCHK, CDN_CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_SI_SDFCHK, CDN_nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_SI_SDFCHK, CDN_nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_nSI_SDFCHK, CDN_nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_SI_SDFCHK, CDN_nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_nSI_SDFCHK, CDN_nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_nSI_SDFCHK, CDN_nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_SI_SDFCHK, CDN_nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_nSI_SDFCHK, CDN_nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_SI_SDFCHK, CDN_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_nSI_SDFCHK, CDN_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SI_SDFCHK, CDN_nD_SDN_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSI_SDFCHK, CDN_D_SDN_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SDFCHK, CDN_D_SDN_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SDFCHK, CDN_nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SDN_SE_SI, CP, D, SDN, SE, SI);
    and (CP_D_SDN_SE_nSI, CP, D, SDN, SE, nSI);
    and (CP_D_SDN_nSE_SI, CP, D, SDN, nSE, SI);
    and (CP_D_SDN_nSE_nSI, CP, D, SDN, nSE, nSI);
    and (CP_nD_SDN_SE_SI, CP, nD, SDN, SE, SI);
    and (CP_nD_SDN_SE_nSI, CP, nD, SDN, SE, nSI);
    and (CP_nD_SDN_nSE_SI, CP, nD, SDN, nSE, SI);
    and (CP_nD_SDN_nSE_nSI, CP, nD, SDN, nSE, nSI);
    and (nCP_D_SDN_SE_SI, nCP, D, SDN, SE, SI);
    and (nCP_D_SDN_SE_nSI, nCP, D, SDN, SE, nSI);
    and (nCP_D_SDN_nSE_SI, nCP, D, SDN, nSE, SI);
    and (nCP_D_SDN_nSE_nSI, nCP, D, SDN, nSE, nSI);
    and (nCP_nD_SDN_SE_SI, nCP, nD, SDN, SE, SI);
    and (nCP_nD_SDN_SE_nSI, nCP, nD, SDN, SE, nSI);
    and (nCP_nD_SDN_nSE_SI, nCP, nD, SDN, nSE, SI);
    and (nCP_nD_SDN_nSE_nSI, nCP, nD, SDN, nSE, nSI);
    and (CDN_D_SDN_SE_SI, CDN, D, SDN, SE, SI);
    and (CDN_D_SDN_nSE_SI, CDN, D, SDN, nSE, SI);
    and (CDN_D_SDN_nSE_nSI, CDN, D, SDN, nSE, nSI);
    and (CDN_nD_SDN_SE_SI, CDN, nD, SDN, SE, SI);
    and (CDN_D_SDN_SE_nSI, CDN, D, SDN, SE, nSI);
    and (CDN_nD_SDN_SE_nSI, CDN, nD, SDN, SE, nSI);
    and (CDN_nD_SDN_nSE_SI, CDN, nD, SDN, nSE, SI);
    and (CDN_nD_SDN_nSE_nSI, CDN, nD, SDN, nSE, nSI);
    and (CDN_CP_D_SE_SI, CDN, CP, D, SE, SI);
    and (CDN_CP_D_SE_nSI, CDN, CP, D, SE, nSI);
    and (CDN_CP_D_nSE_SI, CDN, CP, D, nSE, SI);
    and (CDN_CP_D_nSE_nSI, CDN, CP, D, nSE, nSI);
    and (CDN_CP_nD_SE_SI, CDN, CP, nD, SE, SI);
    and (CDN_CP_nD_SE_nSI, CDN, CP, nD, SE, nSI);
    and (CDN_CP_nD_nSE_SI, CDN, CP, nD, nSE, SI);
    and (CDN_CP_nD_nSE_nSI, CDN, CP, nD, nSE, nSI);
    and (CDN_nCP_D_SE_SI, CDN, nCP, D, SE, SI);
    and (CDN_nCP_D_nSE_SI, CDN, nCP, D, nSE, SI);
    and (CDN_nCP_D_nSE_nSI, CDN, nCP, D, nSE, nSI);
    and (CDN_nCP_nD_SE_SI, CDN, nCP, nD, SE, SI);
    and (CDN_nCP_D_SE_nSI, CDN, nCP, D, SE, nSI);
    and (CDN_nCP_nD_SE_nSI, CDN, nCP, nD, SE, nSI);
    and (CDN_nCP_nD_nSE_SI, CDN, nCP, nD, nSE, SI);
    and (CDN_nCP_nD_nSE_nSI, CDN, nCP, nD, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_SDN_nSE_SI, CDN, SDN, nSE, SI);
    and (CDN_SDN_nSE_nSI, CDN, SDN, nSE, nSI);
    and (CDN_nD_SDN_SI, CDN, nD, SDN, SI);
    and (CDN_D_SDN_nSI, CDN, D, SDN, nSI);
    and (CDN_D_SDN_SE, CDN, D, SDN, SE);
    and (CDN_nD_SDN_SE, CDN, nD, SDN, SE);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SDN_i, SE);
  `endif
  and  (D_check, CDN_i, SDN_i, SE_int_not);
  and  (CP_check, CDN_i, SDN_i);
  and  (SE_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCSNQD4 (SI, D, SE, CP, CDN, SDN, Q);
    input SI, D, SE, CP, CDN, SDN;
    output Q;
    reg notifier;
    reg flag;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SDN_SE_SI_SDFCHK, CP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_SE_nSI_SDFCHK, CP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_SI_SDFCHK, CP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_nSI_SDFCHK, CP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_SI_SDFCHK, CP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_nSI_SDFCHK, CP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_SI_SDFCHK, CP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_nSI_SDFCHK, CP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_SI_SDFCHK, nCP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_nSI_SDFCHK, nCP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_SI_SDFCHK, nCP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_nSI_SDFCHK, nCP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_SI_SDFCHK, nCP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_nSI_SDFCHK, nCP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_SI_SDFCHK, nCP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_nSI_SDFCHK, nCP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SI_SDFCHK, CDN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_SI_SDFCHK, CDN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_nSI_SDFCHK, CDN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SI_SDFCHK, CDN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_nSI_SDFCHK, CDN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_nSI_SDFCHK, CDN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_SI_SDFCHK, CDN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_nSI_SDFCHK, CDN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_SI_SDFCHK, CDN_CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_nSI_SDFCHK, CDN_CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_SI_SDFCHK, CDN_CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_nSI_SDFCHK, CDN_CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_SI_SDFCHK, CDN_CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_nSI_SDFCHK, CDN_CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_SI_SDFCHK, CDN_CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_nSI_SDFCHK, CDN_CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_SI_SDFCHK, CDN_nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_SI_SDFCHK, CDN_nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_nSI_SDFCHK, CDN_nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_SI_SDFCHK, CDN_nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_nSI_SDFCHK, CDN_nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_nSI_SDFCHK, CDN_nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_SI_SDFCHK, CDN_nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_nSI_SDFCHK, CDN_nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_SI_SDFCHK, CDN_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_nSI_SDFCHK, CDN_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SI_SDFCHK, CDN_nD_SDN_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSI_SDFCHK, CDN_D_SDN_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SDFCHK, CDN_D_SDN_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SDFCHK, CDN_nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SDN_SE_SI, CP, D, SDN, SE, SI);
    and (CP_D_SDN_SE_nSI, CP, D, SDN, SE, nSI);
    and (CP_D_SDN_nSE_SI, CP, D, SDN, nSE, SI);
    and (CP_D_SDN_nSE_nSI, CP, D, SDN, nSE, nSI);
    and (CP_nD_SDN_SE_SI, CP, nD, SDN, SE, SI);
    and (CP_nD_SDN_SE_nSI, CP, nD, SDN, SE, nSI);
    and (CP_nD_SDN_nSE_SI, CP, nD, SDN, nSE, SI);
    and (CP_nD_SDN_nSE_nSI, CP, nD, SDN, nSE, nSI);
    and (nCP_D_SDN_SE_SI, nCP, D, SDN, SE, SI);
    and (nCP_D_SDN_SE_nSI, nCP, D, SDN, SE, nSI);
    and (nCP_D_SDN_nSE_SI, nCP, D, SDN, nSE, SI);
    and (nCP_D_SDN_nSE_nSI, nCP, D, SDN, nSE, nSI);
    and (nCP_nD_SDN_SE_SI, nCP, nD, SDN, SE, SI);
    and (nCP_nD_SDN_SE_nSI, nCP, nD, SDN, SE, nSI);
    and (nCP_nD_SDN_nSE_SI, nCP, nD, SDN, nSE, SI);
    and (nCP_nD_SDN_nSE_nSI, nCP, nD, SDN, nSE, nSI);
    and (CDN_D_SDN_SE_SI, CDN, D, SDN, SE, SI);
    and (CDN_D_SDN_nSE_SI, CDN, D, SDN, nSE, SI);
    and (CDN_D_SDN_nSE_nSI, CDN, D, SDN, nSE, nSI);
    and (CDN_nD_SDN_SE_SI, CDN, nD, SDN, SE, SI);
    and (CDN_D_SDN_SE_nSI, CDN, D, SDN, SE, nSI);
    and (CDN_nD_SDN_SE_nSI, CDN, nD, SDN, SE, nSI);
    and (CDN_nD_SDN_nSE_SI, CDN, nD, SDN, nSE, SI);
    and (CDN_nD_SDN_nSE_nSI, CDN, nD, SDN, nSE, nSI);
    and (CDN_CP_D_SE_SI, CDN, CP, D, SE, SI);
    and (CDN_CP_D_SE_nSI, CDN, CP, D, SE, nSI);
    and (CDN_CP_D_nSE_SI, CDN, CP, D, nSE, SI);
    and (CDN_CP_D_nSE_nSI, CDN, CP, D, nSE, nSI);
    and (CDN_CP_nD_SE_SI, CDN, CP, nD, SE, SI);
    and (CDN_CP_nD_SE_nSI, CDN, CP, nD, SE, nSI);
    and (CDN_CP_nD_nSE_SI, CDN, CP, nD, nSE, SI);
    and (CDN_CP_nD_nSE_nSI, CDN, CP, nD, nSE, nSI);
    and (CDN_nCP_D_SE_SI, CDN, nCP, D, SE, SI);
    and (CDN_nCP_D_nSE_SI, CDN, nCP, D, nSE, SI);
    and (CDN_nCP_D_nSE_nSI, CDN, nCP, D, nSE, nSI);
    and (CDN_nCP_nD_SE_SI, CDN, nCP, nD, SE, SI);
    and (CDN_nCP_D_SE_nSI, CDN, nCP, D, SE, nSI);
    and (CDN_nCP_nD_SE_nSI, CDN, nCP, nD, SE, nSI);
    and (CDN_nCP_nD_nSE_SI, CDN, nCP, nD, nSE, SI);
    and (CDN_nCP_nD_nSE_nSI, CDN, nCP, nD, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_SDN_nSE_SI, CDN, SDN, nSE, SI);
    and (CDN_SDN_nSE_nSI, CDN, SDN, nSE, nSI);
    and (CDN_nD_SDN_SI, CDN, nD, SDN, SI);
    and (CDN_D_SDN_nSI, CDN, D, SDN, nSI);
    and (CDN_D_SDN_SE, CDN, D, SDN, SE);
    and (CDN_nD_SDN_SE, CDN, nD, SDN, SE);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SDN_i, SE);
  `endif
  and  (D_check, CDN_i, SDN_i, SE_int_not);
  and  (CP_check, CDN_i, SDN_i);
  and  (SE_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFD0 (SI, D, SE, CP, Q, QN);
    input SI, D, SE, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CP_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFD1 (SI, D, SE, CP, Q, QN);
    input SI, D, SE, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CP_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFD2 (SI, D, SE, CP, Q, QN);
    input SI, D, SE, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CP_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFD4 (SI, D, SE, CP, Q, QN);
    input SI, D, SE, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CP_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCND0 (SI, D, SE, CP, CN, Q, QN);
    input SI, D, SE, CP, CN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        and (D1, CN_d, D_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        and (D1, CN, D);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SE_SI_SDFCHK, CN_D_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SDFCHK, CN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SDFCHK, CN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_SDFCHK, CN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_SDFCHK, nCN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_SDFCHK, nCN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_SDFCHK, CN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_SDFCHK, CN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_SDFCHK, nCN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_SDFCHK, nCN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_SDFCHK, nCN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_SDFCHK, nCN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_SDFCHK, nCN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_SDFCHK, nCN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nSE_SI_SDFCHK, CN_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nSE_nSI_SDFCHK, CN_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SI_SDFCHK, CN_nD_SI, 1'b1);
    tsmc_xbuf (nCN_D_SI_SDFCHK, nCN_D_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SI_SDFCHK, nCN_nD_SI, 1'b1);
    tsmc_xbuf (CN_D_nSI_SDFCHK, CN_D_nSI, 1'b1);
    tsmc_xbuf (CN_D_SE_SDFCHK, CN_D_SE, 1'b1);
    tsmc_xbuf (CN_nD_SE_SDFCHK, CN_nD_SE, 1'b1);
    tsmc_xbuf (nCN_D_SE_SDFCHK, nCN_D_SE, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SDFCHK, nCN_nD_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    and (CN_D_SE_SI, CN, D, SE, SI);
    and (CN_D_nSE_SI, CN, D, nSE, SI);
    and (CN_D_nSE_nSI, CN, D, nSE, nSI);
    and (CN_nD_SE_SI, CN, nD, SE, SI);
    and (nCN_D_SE_SI, nCN, D, SE, SI);
    and (nCN_nD_SE_SI, nCN, nD, SE, SI);
    and (CN_D_SE_nSI, CN, D, SE, nSI);
    and (CN_nD_SE_nSI, CN, nD, SE, nSI);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);
    and (nCN_D_SE_nSI, nCN, D, SE, nSI);
    and (nCN_D_nSE_SI, nCN, D, nSE, SI);
    and (nCN_D_nSE_nSI, nCN, D, nSE, nSI);
    and (nCN_nD_SE_nSI, nCN, nD, SE, nSI);
    and (nCN_nD_nSE_SI, nCN, nD, nSE, SI);
    and (nCN_nD_nSE_nSI, nCN, nD, nSE, nSI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (CN_nSE_SI, CN, nSE, SI);
    and (CN_nSE_nSI, CN, nSE, nSI);
    and (CN_nD_SI, CN, nD, SI);
    and (nCN_D_SI, nCN, D, SI);
    and (nCN_nD_SI, nCN, nD, SI);
    and (CN_D_nSI, CN, D, nSI);
    and (CN_D_SE, CN, D, SE);
    and (CN_nD_SE, CN, nD, SE);
    and (nCN_D_SE, nCN, D, SE);
    and (nCN_nD_SE, nCN, nD, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, CN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, CN);
  `endif
  buf  (CN_check, SE_int_not);
   `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    $width (posedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCND1 (SI, D, SE, CP, CN, Q, QN);
    input SI, D, SE, CP, CN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        and (D1, CN_d, D_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        and (D1, CN, D);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SE_SI_SDFCHK, CN_D_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SDFCHK, CN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SDFCHK, CN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_SDFCHK, CN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_SDFCHK, nCN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_SDFCHK, nCN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_SDFCHK, CN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_SDFCHK, CN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_SDFCHK, nCN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_SDFCHK, nCN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_SDFCHK, nCN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_SDFCHK, nCN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_SDFCHK, nCN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_SDFCHK, nCN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nSE_SI_SDFCHK, CN_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nSE_nSI_SDFCHK, CN_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SI_SDFCHK, CN_nD_SI, 1'b1);
    tsmc_xbuf (nCN_D_SI_SDFCHK, nCN_D_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SI_SDFCHK, nCN_nD_SI, 1'b1);
    tsmc_xbuf (CN_D_nSI_SDFCHK, CN_D_nSI, 1'b1);
    tsmc_xbuf (CN_D_SE_SDFCHK, CN_D_SE, 1'b1);
    tsmc_xbuf (CN_nD_SE_SDFCHK, CN_nD_SE, 1'b1);
    tsmc_xbuf (nCN_D_SE_SDFCHK, nCN_D_SE, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SDFCHK, nCN_nD_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    and (CN_D_SE_SI, CN, D, SE, SI);
    and (CN_D_nSE_SI, CN, D, nSE, SI);
    and (CN_D_nSE_nSI, CN, D, nSE, nSI);
    and (CN_nD_SE_SI, CN, nD, SE, SI);
    and (nCN_D_SE_SI, nCN, D, SE, SI);
    and (nCN_nD_SE_SI, nCN, nD, SE, SI);
    and (CN_D_SE_nSI, CN, D, SE, nSI);
    and (CN_nD_SE_nSI, CN, nD, SE, nSI);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);
    and (nCN_D_SE_nSI, nCN, D, SE, nSI);
    and (nCN_D_nSE_SI, nCN, D, nSE, SI);
    and (nCN_D_nSE_nSI, nCN, D, nSE, nSI);
    and (nCN_nD_SE_nSI, nCN, nD, SE, nSI);
    and (nCN_nD_nSE_SI, nCN, nD, nSE, SI);
    and (nCN_nD_nSE_nSI, nCN, nD, nSE, nSI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (CN_nSE_SI, CN, nSE, SI);
    and (CN_nSE_nSI, CN, nSE, nSI);
    and (CN_nD_SI, CN, nD, SI);
    and (nCN_D_SI, nCN, D, SI);
    and (nCN_nD_SI, nCN, nD, SI);
    and (CN_D_nSI, CN, D, nSI);
    and (CN_D_SE, CN, D, SE);
    and (CN_nD_SE, CN, nD, SE);
    and (nCN_D_SE, nCN, D, SE);
    and (nCN_nD_SE, nCN, nD, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, CN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, CN);
  `endif
  buf  (CN_check, SE_int_not);
   `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    $width (posedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCND2 (SI, D, SE, CP, CN, Q, QN);
    input SI, D, SE, CP, CN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        and (D1, CN_d, D_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        and (D1, CN, D);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SE_SI_SDFCHK, CN_D_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SDFCHK, CN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SDFCHK, CN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_SDFCHK, CN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_SDFCHK, nCN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_SDFCHK, nCN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_SDFCHK, CN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_SDFCHK, CN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_SDFCHK, nCN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_SDFCHK, nCN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_SDFCHK, nCN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_SDFCHK, nCN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_SDFCHK, nCN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_SDFCHK, nCN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nSE_SI_SDFCHK, CN_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nSE_nSI_SDFCHK, CN_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SI_SDFCHK, CN_nD_SI, 1'b1);
    tsmc_xbuf (nCN_D_SI_SDFCHK, nCN_D_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SI_SDFCHK, nCN_nD_SI, 1'b1);
    tsmc_xbuf (CN_D_nSI_SDFCHK, CN_D_nSI, 1'b1);
    tsmc_xbuf (CN_D_SE_SDFCHK, CN_D_SE, 1'b1);
    tsmc_xbuf (CN_nD_SE_SDFCHK, CN_nD_SE, 1'b1);
    tsmc_xbuf (nCN_D_SE_SDFCHK, nCN_D_SE, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SDFCHK, nCN_nD_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    and (CN_D_SE_SI, CN, D, SE, SI);
    and (CN_D_nSE_SI, CN, D, nSE, SI);
    and (CN_D_nSE_nSI, CN, D, nSE, nSI);
    and (CN_nD_SE_SI, CN, nD, SE, SI);
    and (nCN_D_SE_SI, nCN, D, SE, SI);
    and (nCN_nD_SE_SI, nCN, nD, SE, SI);
    and (CN_D_SE_nSI, CN, D, SE, nSI);
    and (CN_nD_SE_nSI, CN, nD, SE, nSI);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);
    and (nCN_D_SE_nSI, nCN, D, SE, nSI);
    and (nCN_D_nSE_SI, nCN, D, nSE, SI);
    and (nCN_D_nSE_nSI, nCN, D, nSE, nSI);
    and (nCN_nD_SE_nSI, nCN, nD, SE, nSI);
    and (nCN_nD_nSE_SI, nCN, nD, nSE, SI);
    and (nCN_nD_nSE_nSI, nCN, nD, nSE, nSI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (CN_nSE_SI, CN, nSE, SI);
    and (CN_nSE_nSI, CN, nSE, nSI);
    and (CN_nD_SI, CN, nD, SI);
    and (nCN_D_SI, nCN, D, SI);
    and (nCN_nD_SI, nCN, nD, SI);
    and (CN_D_nSI, CN, D, nSI);
    and (CN_D_SE, CN, D, SE);
    and (CN_nD_SE, CN, nD, SE);
    and (nCN_D_SE, nCN, D, SE);
    and (nCN_nD_SE, nCN, nD, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, CN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, CN);
  `endif
  buf  (CN_check, SE_int_not);
   `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    $width (posedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCND4 (SI, D, SE, CP, CN, Q, QN);
    input SI, D, SE, CP, CN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        and (D1, CN_d, D_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        and (D1, CN, D);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SE_SI_SDFCHK, CN_D_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SDFCHK, CN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SDFCHK, CN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_SDFCHK, CN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_SDFCHK, nCN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_SDFCHK, nCN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_SDFCHK, CN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_SDFCHK, CN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_SDFCHK, nCN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_SDFCHK, nCN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_SDFCHK, nCN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_SDFCHK, nCN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_SDFCHK, nCN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_SDFCHK, nCN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nSE_SI_SDFCHK, CN_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nSE_nSI_SDFCHK, CN_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SI_SDFCHK, CN_nD_SI, 1'b1);
    tsmc_xbuf (nCN_D_SI_SDFCHK, nCN_D_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SI_SDFCHK, nCN_nD_SI, 1'b1);
    tsmc_xbuf (CN_D_nSI_SDFCHK, CN_D_nSI, 1'b1);
    tsmc_xbuf (CN_D_SE_SDFCHK, CN_D_SE, 1'b1);
    tsmc_xbuf (CN_nD_SE_SDFCHK, CN_nD_SE, 1'b1);
    tsmc_xbuf (nCN_D_SE_SDFCHK, nCN_D_SE, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SDFCHK, nCN_nD_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    and (CN_D_SE_SI, CN, D, SE, SI);
    and (CN_D_nSE_SI, CN, D, nSE, SI);
    and (CN_D_nSE_nSI, CN, D, nSE, nSI);
    and (CN_nD_SE_SI, CN, nD, SE, SI);
    and (nCN_D_SE_SI, nCN, D, SE, SI);
    and (nCN_nD_SE_SI, nCN, nD, SE, SI);
    and (CN_D_SE_nSI, CN, D, SE, nSI);
    and (CN_nD_SE_nSI, CN, nD, SE, nSI);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);
    and (nCN_D_SE_nSI, nCN, D, SE, nSI);
    and (nCN_D_nSE_SI, nCN, D, nSE, SI);
    and (nCN_D_nSE_nSI, nCN, D, nSE, nSI);
    and (nCN_nD_SE_nSI, nCN, nD, SE, nSI);
    and (nCN_nD_nSE_SI, nCN, nD, nSE, SI);
    and (nCN_nD_nSE_nSI, nCN, nD, nSE, nSI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (CN_nSE_SI, CN, nSE, SI);
    and (CN_nSE_nSI, CN, nSE, nSI);
    and (CN_nD_SI, CN, nD, SI);
    and (nCN_D_SI, nCN, D, SI);
    and (nCN_nD_SI, nCN, nD, SI);
    and (CN_D_nSI, CN, D, nSI);
    and (CN_D_SE, CN, D, SE);
    and (CN_nD_SE, CN, nD, SE);
    and (nCN_D_SE, nCN, D, SE);
    and (nCN_nD_SE, nCN, nD, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, CN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, CN);
  `endif
  buf  (CN_check, SE_int_not);
   `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    $width (posedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCNQD0 (SI, D, SE, CP, CN, Q);
    input SI, D, SE, CP, CN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        and (D1, CN_d, D_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        and (D1, CN, D);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SE_SI_SDFCHK, CN_D_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SDFCHK, CN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SDFCHK, CN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_SDFCHK, CN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_SDFCHK, nCN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_SDFCHK, nCN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_SDFCHK, CN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_SDFCHK, CN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_SDFCHK, nCN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_SDFCHK, nCN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_SDFCHK, nCN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_SDFCHK, nCN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_SDFCHK, nCN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_SDFCHK, nCN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nSE_SI_SDFCHK, CN_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nSE_nSI_SDFCHK, CN_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SI_SDFCHK, CN_nD_SI, 1'b1);
    tsmc_xbuf (nCN_D_SI_SDFCHK, nCN_D_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SI_SDFCHK, nCN_nD_SI, 1'b1);
    tsmc_xbuf (CN_D_nSI_SDFCHK, CN_D_nSI, 1'b1);
    tsmc_xbuf (CN_D_SE_SDFCHK, CN_D_SE, 1'b1);
    tsmc_xbuf (CN_nD_SE_SDFCHK, CN_nD_SE, 1'b1);
    tsmc_xbuf (nCN_D_SE_SDFCHK, nCN_D_SE, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SDFCHK, nCN_nD_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    and (CN_D_SE_SI, CN, D, SE, SI);
    and (CN_D_nSE_SI, CN, D, nSE, SI);
    and (CN_D_nSE_nSI, CN, D, nSE, nSI);
    and (CN_nD_SE_SI, CN, nD, SE, SI);
    and (nCN_D_SE_SI, nCN, D, SE, SI);
    and (nCN_nD_SE_SI, nCN, nD, SE, SI);
    and (CN_D_SE_nSI, CN, D, SE, nSI);
    and (CN_nD_SE_nSI, CN, nD, SE, nSI);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);
    and (nCN_D_SE_nSI, nCN, D, SE, nSI);
    and (nCN_D_nSE_SI, nCN, D, nSE, SI);
    and (nCN_D_nSE_nSI, nCN, D, nSE, nSI);
    and (nCN_nD_SE_nSI, nCN, nD, SE, nSI);
    and (nCN_nD_nSE_SI, nCN, nD, nSE, SI);
    and (nCN_nD_nSE_nSI, nCN, nD, nSE, nSI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (CN_nSE_SI, CN, nSE, SI);
    and (CN_nSE_nSI, CN, nSE, nSI);
    and (CN_nD_SI, CN, nD, SI);
    and (nCN_D_SI, nCN, D, SI);
    and (nCN_nD_SI, nCN, nD, SI);
    and (CN_D_nSI, CN, D, nSI);
    and (CN_D_SE, CN, D, SE);
    and (CN_nD_SE, CN, nD, SE);
    and (nCN_D_SE, nCN, D, SE);
    and (nCN_nD_SE, nCN, nD, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, CN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, CN);
  `endif
  buf  (CN_check, SE_int_not);
   `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    $width (posedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCNQD1 (SI, D, SE, CP, CN, Q);
    input SI, D, SE, CP, CN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        and (D1, CN_d, D_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        and (D1, CN, D);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SE_SI_SDFCHK, CN_D_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SDFCHK, CN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SDFCHK, CN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_SDFCHK, CN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_SDFCHK, nCN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_SDFCHK, nCN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_SDFCHK, CN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_SDFCHK, CN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_SDFCHK, nCN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_SDFCHK, nCN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_SDFCHK, nCN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_SDFCHK, nCN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_SDFCHK, nCN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_SDFCHK, nCN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nSE_SI_SDFCHK, CN_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nSE_nSI_SDFCHK, CN_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SI_SDFCHK, CN_nD_SI, 1'b1);
    tsmc_xbuf (nCN_D_SI_SDFCHK, nCN_D_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SI_SDFCHK, nCN_nD_SI, 1'b1);
    tsmc_xbuf (CN_D_nSI_SDFCHK, CN_D_nSI, 1'b1);
    tsmc_xbuf (CN_D_SE_SDFCHK, CN_D_SE, 1'b1);
    tsmc_xbuf (CN_nD_SE_SDFCHK, CN_nD_SE, 1'b1);
    tsmc_xbuf (nCN_D_SE_SDFCHK, nCN_D_SE, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SDFCHK, nCN_nD_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    and (CN_D_SE_SI, CN, D, SE, SI);
    and (CN_D_nSE_SI, CN, D, nSE, SI);
    and (CN_D_nSE_nSI, CN, D, nSE, nSI);
    and (CN_nD_SE_SI, CN, nD, SE, SI);
    and (nCN_D_SE_SI, nCN, D, SE, SI);
    and (nCN_nD_SE_SI, nCN, nD, SE, SI);
    and (CN_D_SE_nSI, CN, D, SE, nSI);
    and (CN_nD_SE_nSI, CN, nD, SE, nSI);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);
    and (nCN_D_SE_nSI, nCN, D, SE, nSI);
    and (nCN_D_nSE_SI, nCN, D, nSE, SI);
    and (nCN_D_nSE_nSI, nCN, D, nSE, nSI);
    and (nCN_nD_SE_nSI, nCN, nD, SE, nSI);
    and (nCN_nD_nSE_SI, nCN, nD, nSE, SI);
    and (nCN_nD_nSE_nSI, nCN, nD, nSE, nSI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (CN_nSE_SI, CN, nSE, SI);
    and (CN_nSE_nSI, CN, nSE, nSI);
    and (CN_nD_SI, CN, nD, SI);
    and (nCN_D_SI, nCN, D, SI);
    and (nCN_nD_SI, nCN, nD, SI);
    and (CN_D_nSI, CN, D, nSI);
    and (CN_D_SE, CN, D, SE);
    and (CN_nD_SE, CN, nD, SE);
    and (nCN_D_SE, nCN, D, SE);
    and (nCN_nD_SE, nCN, nD, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, CN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, CN);
  `endif
  buf  (CN_check, SE_int_not);
   `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    $width (posedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCNQD2 (SI, D, SE, CP, CN, Q);
    input SI, D, SE, CP, CN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        and (D1, CN_d, D_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        and (D1, CN, D);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SE_SI_SDFCHK, CN_D_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SDFCHK, CN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SDFCHK, CN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_SDFCHK, CN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_SDFCHK, nCN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_SDFCHK, nCN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_SDFCHK, CN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_SDFCHK, CN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_SDFCHK, nCN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_SDFCHK, nCN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_SDFCHK, nCN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_SDFCHK, nCN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_SDFCHK, nCN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_SDFCHK, nCN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nSE_SI_SDFCHK, CN_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nSE_nSI_SDFCHK, CN_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SI_SDFCHK, CN_nD_SI, 1'b1);
    tsmc_xbuf (nCN_D_SI_SDFCHK, nCN_D_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SI_SDFCHK, nCN_nD_SI, 1'b1);
    tsmc_xbuf (CN_D_nSI_SDFCHK, CN_D_nSI, 1'b1);
    tsmc_xbuf (CN_D_SE_SDFCHK, CN_D_SE, 1'b1);
    tsmc_xbuf (CN_nD_SE_SDFCHK, CN_nD_SE, 1'b1);
    tsmc_xbuf (nCN_D_SE_SDFCHK, nCN_D_SE, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SDFCHK, nCN_nD_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    and (CN_D_SE_SI, CN, D, SE, SI);
    and (CN_D_nSE_SI, CN, D, nSE, SI);
    and (CN_D_nSE_nSI, CN, D, nSE, nSI);
    and (CN_nD_SE_SI, CN, nD, SE, SI);
    and (nCN_D_SE_SI, nCN, D, SE, SI);
    and (nCN_nD_SE_SI, nCN, nD, SE, SI);
    and (CN_D_SE_nSI, CN, D, SE, nSI);
    and (CN_nD_SE_nSI, CN, nD, SE, nSI);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);
    and (nCN_D_SE_nSI, nCN, D, SE, nSI);
    and (nCN_D_nSE_SI, nCN, D, nSE, SI);
    and (nCN_D_nSE_nSI, nCN, D, nSE, nSI);
    and (nCN_nD_SE_nSI, nCN, nD, SE, nSI);
    and (nCN_nD_nSE_SI, nCN, nD, nSE, SI);
    and (nCN_nD_nSE_nSI, nCN, nD, nSE, nSI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (CN_nSE_SI, CN, nSE, SI);
    and (CN_nSE_nSI, CN, nSE, nSI);
    and (CN_nD_SI, CN, nD, SI);
    and (nCN_D_SI, nCN, D, SI);
    and (nCN_nD_SI, nCN, nD, SI);
    and (CN_D_nSI, CN, D, nSI);
    and (CN_D_SE, CN, D, SE);
    and (CN_nD_SE, CN, nD, SE);
    and (nCN_D_SE, nCN, D, SE);
    and (nCN_nD_SE, nCN, nD, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, CN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, CN);
  `endif
  buf  (CN_check, SE_int_not);
   `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    $width (posedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCNQD4 (SI, D, SE, CP, CN, Q);
    input SI, D, SE, CP, CN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        and (D1, CN_d, D_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        and (D1, CN, D);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SE_SI_SDFCHK, CN_D_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SDFCHK, CN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SDFCHK, CN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_SDFCHK, CN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_SDFCHK, nCN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_SDFCHK, nCN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_SDFCHK, CN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_SDFCHK, CN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_SDFCHK, nCN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_SDFCHK, nCN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_SDFCHK, nCN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_SDFCHK, nCN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_SDFCHK, nCN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_SDFCHK, nCN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nSE_SI_SDFCHK, CN_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nSE_nSI_SDFCHK, CN_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SI_SDFCHK, CN_nD_SI, 1'b1);
    tsmc_xbuf (nCN_D_SI_SDFCHK, nCN_D_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SI_SDFCHK, nCN_nD_SI, 1'b1);
    tsmc_xbuf (CN_D_nSI_SDFCHK, CN_D_nSI, 1'b1);
    tsmc_xbuf (CN_D_SE_SDFCHK, CN_D_SE, 1'b1);
    tsmc_xbuf (CN_nD_SE_SDFCHK, CN_nD_SE, 1'b1);
    tsmc_xbuf (nCN_D_SE_SDFCHK, nCN_D_SE, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SDFCHK, nCN_nD_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    and (CN_D_SE_SI, CN, D, SE, SI);
    and (CN_D_nSE_SI, CN, D, nSE, SI);
    and (CN_D_nSE_nSI, CN, D, nSE, nSI);
    and (CN_nD_SE_SI, CN, nD, SE, SI);
    and (nCN_D_SE_SI, nCN, D, SE, SI);
    and (nCN_nD_SE_SI, nCN, nD, SE, SI);
    and (CN_D_SE_nSI, CN, D, SE, nSI);
    and (CN_nD_SE_nSI, CN, nD, SE, nSI);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);
    and (nCN_D_SE_nSI, nCN, D, SE, nSI);
    and (nCN_D_nSE_SI, nCN, D, nSE, SI);
    and (nCN_D_nSE_nSI, nCN, D, nSE, nSI);
    and (nCN_nD_SE_nSI, nCN, nD, SE, nSI);
    and (nCN_nD_nSE_SI, nCN, nD, nSE, SI);
    and (nCN_nD_nSE_nSI, nCN, nD, nSE, nSI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (CN_nSE_SI, CN, nSE, SI);
    and (CN_nSE_nSI, CN, nSE, nSI);
    and (CN_nD_SI, CN, nD, SI);
    and (nCN_D_SI, nCN, D, SI);
    and (nCN_nD_SI, nCN, nD, SI);
    and (CN_D_nSI, CN, D, nSI);
    and (CN_D_SE, CN, D, SE);
    and (CN_nD_SE, CN, nD, SE);
    and (nCN_D_SE, nCN, D, SE);
    and (nCN_nD_SE, nCN, nD, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, CN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, CN);
  `endif
  buf  (CN_check, SE_int_not);
   `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    $width (posedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCSND0 (SI, D, SE, CP, CN, SN, Q, QN);
    input SI, D, SE, CP, CN, SN;
    output Q, QN;
    reg notifier;
    reg flag;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (DS, S, D_d);
        and (D1, DS, CN_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (DS, S, D);
        and (D1, DS, CN);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 
    buf (CN_i, CN);
    buf (SN_i, SN);
    always @(CN_i or SN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CN_i===1'b0)&&(SN_i===1'b0));
            if (flag == 1) begin 
                if (CN_i!==1'b0) begin
                    $display("%m > CN is released at time %.2fns.", $realtime);
                end 
                if (SN_i!==1'b0) begin
                    $display("%m > SN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CN and SN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SE_SI_SN_SDFCHK, CN_D_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_SI_nSN_SDFCHK, CN_D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SN_SDFCHK, CN_D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_nSN_SDFCHK, CN_D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SN_SDFCHK, CN_D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_nSN_SDFCHK, CN_D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_SN_SDFCHK, CN_nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_nSN_SDFCHK, CN_nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_nSN_SDFCHK, CN_nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_nSN_SDFCHK, CN_nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_SN_SDFCHK, nCN_D_SE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_SN_SDFCHK, nCN_nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_SN_SDFCHK, CN_D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_nSN_SDFCHK, CN_D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_SN_SDFCHK, CN_nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_nSN_SDFCHK, CN_nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SN_SDFCHK, CN_nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SN_SDFCHK, CN_nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_SN_SDFCHK, nCN_D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_SN_SDFCHK, nCN_D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_SN_SDFCHK, nCN_D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_SN_SDFCHK, nCN_nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_SN_SDFCHK, nCN_nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_SN_SDFCHK, nCN_nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSE_SI_SN_SDFCHK, D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SN_SDFCHK, D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nSE_SI_SN_SDFCHK, CN_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nSE_nSI_SN_SDFCHK, CN_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SI_SN_SDFCHK, CN_nD_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SI_SN_SDFCHK, nCN_D_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SI_SN_SDFCHK, nCN_nD_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSI_SN_SDFCHK, CN_D_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSI_nSN_SDFCHK, CN_D_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSI_nSN_SDFCHK, CN_nD_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_D_SE_SN_SDFCHK, CN_D_SE_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSN_SDFCHK, CN_D_SE_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SN_SDFCHK, CN_nD_SE_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSN_SDFCHK, CN_nD_SE_nSN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SN_SDFCHK, nCN_D_SE_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SN_SDFCHK, nCN_nD_SE_SN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    not (nSN, SN);
    and (CN_D_SE_SI_SN, CN, D, SE, SI, SN);
    and (CN_D_SE_SI_nSN, CN, D, SE, SI, nSN);
    and (CN_D_nSE_SI_SN, CN, D, nSE, SI, SN);
    and (CN_D_nSE_SI_nSN, CN, D, nSE, SI, nSN);
    and (CN_D_nSE_nSI_SN, CN, D, nSE, nSI, SN);
    and (CN_D_nSE_nSI_nSN, CN, D, nSE, nSI, nSN);
    and (CN_nD_SE_SI_SN, CN, nD, SE, SI, SN);
    and (CN_nD_SE_SI_nSN, CN, nD, SE, SI, nSN);
    and (CN_nD_nSE_SI_nSN, CN, nD, nSE, SI, nSN);
    and (CN_nD_nSE_nSI_nSN, CN, nD, nSE, nSI, nSN);
    and (nCN_D_SE_SI_SN, nCN, D, SE, SI, SN);
    and (nCN_nD_SE_SI_SN, nCN, nD, SE, SI, SN);
    and (CN_D_SE_nSI_SN, CN, D, SE, nSI, SN);
    and (CN_D_SE_nSI_nSN, CN, D, SE, nSI, nSN);
    and (CN_nD_SE_nSI_SN, CN, nD, SE, nSI, SN);
    and (CN_nD_SE_nSI_nSN, CN, nD, SE, nSI, nSN);
    and (CN_nD_nSE_SI_SN, CN, nD, nSE, SI, SN);
    and (CN_nD_nSE_nSI_SN, CN, nD, nSE, nSI, SN);
    and (nCN_D_SE_nSI_SN, nCN, D, SE, nSI, SN);
    and (nCN_D_nSE_SI_SN, nCN, D, nSE, SI, SN);
    and (nCN_D_nSE_nSI_SN, nCN, D, nSE, nSI, SN);
    and (nCN_nD_SE_nSI_SN, nCN, nD, SE, nSI, SN);
    and (nCN_nD_nSE_SI_SN, nCN, nD, nSE, SI, SN);
    and (nCN_nD_nSE_nSI_SN, nCN, nD, nSE, nSI, SN);
    and (D_nSE_SI_SN, D, nSE, SI, SN);
    and (D_nSE_nSI_SN, D, nSE, nSI, SN);
    and (CN_nSE_SI_SN, CN, nSE, SI, SN);
    and (CN_nSE_nSI_SN, CN, nSE, nSI, SN);
    and (CN_nD_SI_SN, CN, nD, SI, SN);
    and (nCN_D_SI_SN, nCN, D, SI, SN);
    and (nCN_nD_SI_SN, nCN, nD, SI, SN);
    and (CN_D_nSI_SN, CN, D, nSI, SN);
    and (CN_D_nSI_nSN, CN, D, nSI, nSN);
    and (CN_nD_nSI_nSN, CN, nD, nSI, nSN);
    and (CN_D_SE_SN, CN, D, SE, SN);
    and (CN_D_SE_nSN, CN, D, SE, nSN);
    and (CN_nD_SE_SN, CN, nD, SE, SN);
    and (CN_nD_SE_nSN, CN, nD, SE, nSN);
    and (nCN_D_SE_SN, nCN, D, SE, SN);
    and (nCN_nD_SE_SN, nCN, nD, SE, SN);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, CN_d, SN_d);
    and  (SN_check, SE_int_not, CN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, CN, SN);
    and  (SN_check, SE_int_not, CN);
  `endif
  buf  (CN_check, SE_int_not);
   `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& CN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCSND1 (SI, D, SE, CP, CN, SN, Q, QN);
    input SI, D, SE, CP, CN, SN;
    output Q, QN;
    reg notifier;
    reg flag;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (DS, S, D_d);
        and (D1, DS, CN_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (DS, S, D);
        and (D1, DS, CN);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 
    buf (CN_i, CN);
    buf (SN_i, SN);
    always @(CN_i or SN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CN_i===1'b0)&&(SN_i===1'b0));
            if (flag == 1) begin 
                if (CN_i!==1'b0) begin
                    $display("%m > CN is released at time %.2fns.", $realtime);
                end 
                if (SN_i!==1'b0) begin
                    $display("%m > SN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CN and SN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SE_SI_SN_SDFCHK, CN_D_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_SI_nSN_SDFCHK, CN_D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SN_SDFCHK, CN_D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_nSN_SDFCHK, CN_D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SN_SDFCHK, CN_D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_nSN_SDFCHK, CN_D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_SN_SDFCHK, CN_nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_nSN_SDFCHK, CN_nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_nSN_SDFCHK, CN_nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_nSN_SDFCHK, CN_nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_SN_SDFCHK, nCN_D_SE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_SN_SDFCHK, nCN_nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_SN_SDFCHK, CN_D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_nSN_SDFCHK, CN_D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_SN_SDFCHK, CN_nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_nSN_SDFCHK, CN_nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SN_SDFCHK, CN_nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SN_SDFCHK, CN_nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_SN_SDFCHK, nCN_D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_SN_SDFCHK, nCN_D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_SN_SDFCHK, nCN_D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_SN_SDFCHK, nCN_nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_SN_SDFCHK, nCN_nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_SN_SDFCHK, nCN_nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSE_SI_SN_SDFCHK, D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SN_SDFCHK, D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nSE_SI_SN_SDFCHK, CN_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nSE_nSI_SN_SDFCHK, CN_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SI_SN_SDFCHK, CN_nD_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SI_SN_SDFCHK, nCN_D_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SI_SN_SDFCHK, nCN_nD_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSI_SN_SDFCHK, CN_D_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSI_nSN_SDFCHK, CN_D_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSI_nSN_SDFCHK, CN_nD_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_D_SE_SN_SDFCHK, CN_D_SE_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSN_SDFCHK, CN_D_SE_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SN_SDFCHK, CN_nD_SE_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSN_SDFCHK, CN_nD_SE_nSN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SN_SDFCHK, nCN_D_SE_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SN_SDFCHK, nCN_nD_SE_SN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    not (nSN, SN);
    and (CN_D_SE_SI_SN, CN, D, SE, SI, SN);
    and (CN_D_SE_SI_nSN, CN, D, SE, SI, nSN);
    and (CN_D_nSE_SI_SN, CN, D, nSE, SI, SN);
    and (CN_D_nSE_SI_nSN, CN, D, nSE, SI, nSN);
    and (CN_D_nSE_nSI_SN, CN, D, nSE, nSI, SN);
    and (CN_D_nSE_nSI_nSN, CN, D, nSE, nSI, nSN);
    and (CN_nD_SE_SI_SN, CN, nD, SE, SI, SN);
    and (CN_nD_SE_SI_nSN, CN, nD, SE, SI, nSN);
    and (CN_nD_nSE_SI_nSN, CN, nD, nSE, SI, nSN);
    and (CN_nD_nSE_nSI_nSN, CN, nD, nSE, nSI, nSN);
    and (nCN_D_SE_SI_SN, nCN, D, SE, SI, SN);
    and (nCN_nD_SE_SI_SN, nCN, nD, SE, SI, SN);
    and (CN_D_SE_nSI_SN, CN, D, SE, nSI, SN);
    and (CN_D_SE_nSI_nSN, CN, D, SE, nSI, nSN);
    and (CN_nD_SE_nSI_SN, CN, nD, SE, nSI, SN);
    and (CN_nD_SE_nSI_nSN, CN, nD, SE, nSI, nSN);
    and (CN_nD_nSE_SI_SN, CN, nD, nSE, SI, SN);
    and (CN_nD_nSE_nSI_SN, CN, nD, nSE, nSI, SN);
    and (nCN_D_SE_nSI_SN, nCN, D, SE, nSI, SN);
    and (nCN_D_nSE_SI_SN, nCN, D, nSE, SI, SN);
    and (nCN_D_nSE_nSI_SN, nCN, D, nSE, nSI, SN);
    and (nCN_nD_SE_nSI_SN, nCN, nD, SE, nSI, SN);
    and (nCN_nD_nSE_SI_SN, nCN, nD, nSE, SI, SN);
    and (nCN_nD_nSE_nSI_SN, nCN, nD, nSE, nSI, SN);
    and (D_nSE_SI_SN, D, nSE, SI, SN);
    and (D_nSE_nSI_SN, D, nSE, nSI, SN);
    and (CN_nSE_SI_SN, CN, nSE, SI, SN);
    and (CN_nSE_nSI_SN, CN, nSE, nSI, SN);
    and (CN_nD_SI_SN, CN, nD, SI, SN);
    and (nCN_D_SI_SN, nCN, D, SI, SN);
    and (nCN_nD_SI_SN, nCN, nD, SI, SN);
    and (CN_D_nSI_SN, CN, D, nSI, SN);
    and (CN_D_nSI_nSN, CN, D, nSI, nSN);
    and (CN_nD_nSI_nSN, CN, nD, nSI, nSN);
    and (CN_D_SE_SN, CN, D, SE, SN);
    and (CN_D_SE_nSN, CN, D, SE, nSN);
    and (CN_nD_SE_SN, CN, nD, SE, SN);
    and (CN_nD_SE_nSN, CN, nD, SE, nSN);
    and (nCN_D_SE_SN, nCN, D, SE, SN);
    and (nCN_nD_SE_SN, nCN, nD, SE, SN);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, CN_d, SN_d);
    and  (SN_check, SE_int_not, CN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, CN, SN);
    and  (SN_check, SE_int_not, CN);
  `endif
  buf  (CN_check, SE_int_not);
   `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& CN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCSND2 (SI, D, SE, CP, CN, SN, Q, QN);
    input SI, D, SE, CP, CN, SN;
    output Q, QN;
    reg notifier;
    reg flag;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (DS, S, D_d);
        and (D1, DS, CN_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (DS, S, D);
        and (D1, DS, CN);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 
    buf (CN_i, CN);
    buf (SN_i, SN);
    always @(CN_i or SN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CN_i===1'b0)&&(SN_i===1'b0));
            if (flag == 1) begin 
                if (CN_i!==1'b0) begin
                    $display("%m > CN is released at time %.2fns.", $realtime);
                end 
                if (SN_i!==1'b0) begin
                    $display("%m > SN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CN and SN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SE_SI_SN_SDFCHK, CN_D_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_SI_nSN_SDFCHK, CN_D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SN_SDFCHK, CN_D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_nSN_SDFCHK, CN_D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SN_SDFCHK, CN_D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_nSN_SDFCHK, CN_D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_SN_SDFCHK, CN_nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_nSN_SDFCHK, CN_nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_nSN_SDFCHK, CN_nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_nSN_SDFCHK, CN_nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_SN_SDFCHK, nCN_D_SE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_SN_SDFCHK, nCN_nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_SN_SDFCHK, CN_D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_nSN_SDFCHK, CN_D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_SN_SDFCHK, CN_nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_nSN_SDFCHK, CN_nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SN_SDFCHK, CN_nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SN_SDFCHK, CN_nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_SN_SDFCHK, nCN_D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_SN_SDFCHK, nCN_D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_SN_SDFCHK, nCN_D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_SN_SDFCHK, nCN_nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_SN_SDFCHK, nCN_nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_SN_SDFCHK, nCN_nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSE_SI_SN_SDFCHK, D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SN_SDFCHK, D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nSE_SI_SN_SDFCHK, CN_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nSE_nSI_SN_SDFCHK, CN_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SI_SN_SDFCHK, CN_nD_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SI_SN_SDFCHK, nCN_D_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SI_SN_SDFCHK, nCN_nD_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSI_SN_SDFCHK, CN_D_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSI_nSN_SDFCHK, CN_D_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSI_nSN_SDFCHK, CN_nD_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_D_SE_SN_SDFCHK, CN_D_SE_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSN_SDFCHK, CN_D_SE_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SN_SDFCHK, CN_nD_SE_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSN_SDFCHK, CN_nD_SE_nSN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SN_SDFCHK, nCN_D_SE_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SN_SDFCHK, nCN_nD_SE_SN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    not (nSN, SN);
    and (CN_D_SE_SI_SN, CN, D, SE, SI, SN);
    and (CN_D_SE_SI_nSN, CN, D, SE, SI, nSN);
    and (CN_D_nSE_SI_SN, CN, D, nSE, SI, SN);
    and (CN_D_nSE_SI_nSN, CN, D, nSE, SI, nSN);
    and (CN_D_nSE_nSI_SN, CN, D, nSE, nSI, SN);
    and (CN_D_nSE_nSI_nSN, CN, D, nSE, nSI, nSN);
    and (CN_nD_SE_SI_SN, CN, nD, SE, SI, SN);
    and (CN_nD_SE_SI_nSN, CN, nD, SE, SI, nSN);
    and (CN_nD_nSE_SI_nSN, CN, nD, nSE, SI, nSN);
    and (CN_nD_nSE_nSI_nSN, CN, nD, nSE, nSI, nSN);
    and (nCN_D_SE_SI_SN, nCN, D, SE, SI, SN);
    and (nCN_nD_SE_SI_SN, nCN, nD, SE, SI, SN);
    and (CN_D_SE_nSI_SN, CN, D, SE, nSI, SN);
    and (CN_D_SE_nSI_nSN, CN, D, SE, nSI, nSN);
    and (CN_nD_SE_nSI_SN, CN, nD, SE, nSI, SN);
    and (CN_nD_SE_nSI_nSN, CN, nD, SE, nSI, nSN);
    and (CN_nD_nSE_SI_SN, CN, nD, nSE, SI, SN);
    and (CN_nD_nSE_nSI_SN, CN, nD, nSE, nSI, SN);
    and (nCN_D_SE_nSI_SN, nCN, D, SE, nSI, SN);
    and (nCN_D_nSE_SI_SN, nCN, D, nSE, SI, SN);
    and (nCN_D_nSE_nSI_SN, nCN, D, nSE, nSI, SN);
    and (nCN_nD_SE_nSI_SN, nCN, nD, SE, nSI, SN);
    and (nCN_nD_nSE_SI_SN, nCN, nD, nSE, SI, SN);
    and (nCN_nD_nSE_nSI_SN, nCN, nD, nSE, nSI, SN);
    and (D_nSE_SI_SN, D, nSE, SI, SN);
    and (D_nSE_nSI_SN, D, nSE, nSI, SN);
    and (CN_nSE_SI_SN, CN, nSE, SI, SN);
    and (CN_nSE_nSI_SN, CN, nSE, nSI, SN);
    and (CN_nD_SI_SN, CN, nD, SI, SN);
    and (nCN_D_SI_SN, nCN, D, SI, SN);
    and (nCN_nD_SI_SN, nCN, nD, SI, SN);
    and (CN_D_nSI_SN, CN, D, nSI, SN);
    and (CN_D_nSI_nSN, CN, D, nSI, nSN);
    and (CN_nD_nSI_nSN, CN, nD, nSI, nSN);
    and (CN_D_SE_SN, CN, D, SE, SN);
    and (CN_D_SE_nSN, CN, D, SE, nSN);
    and (CN_nD_SE_SN, CN, nD, SE, SN);
    and (CN_nD_SE_nSN, CN, nD, SE, nSN);
    and (nCN_D_SE_SN, nCN, D, SE, SN);
    and (nCN_nD_SE_SN, nCN, nD, SE, SN);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, CN_d, SN_d);
    and  (SN_check, SE_int_not, CN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, CN, SN);
    and  (SN_check, SE_int_not, CN);
  `endif
  buf  (CN_check, SE_int_not);
   `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& CN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCSND4 (SI, D, SE, CP, CN, SN, Q, QN);
    input SI, D, SE, CP, CN, SN;
    output Q, QN;
    reg notifier;
    reg flag;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (DS, S, D_d);
        and (D1, DS, CN_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (DS, S, D);
        and (D1, DS, CN);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 
    buf (CN_i, CN);
    buf (SN_i, SN);
    always @(CN_i or SN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CN_i===1'b0)&&(SN_i===1'b0));
            if (flag == 1) begin 
                if (CN_i!==1'b0) begin
                    $display("%m > CN is released at time %.2fns.", $realtime);
                end 
                if (SN_i!==1'b0) begin
                    $display("%m > SN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CN and SN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SE_SI_SN_SDFCHK, CN_D_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_SI_nSN_SDFCHK, CN_D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SN_SDFCHK, CN_D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_nSN_SDFCHK, CN_D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SN_SDFCHK, CN_D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_nSN_SDFCHK, CN_D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_SN_SDFCHK, CN_nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_nSN_SDFCHK, CN_nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_nSN_SDFCHK, CN_nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_nSN_SDFCHK, CN_nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_SN_SDFCHK, nCN_D_SE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_SN_SDFCHK, nCN_nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_SN_SDFCHK, CN_D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_nSN_SDFCHK, CN_D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_SN_SDFCHK, CN_nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_nSN_SDFCHK, CN_nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SN_SDFCHK, CN_nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SN_SDFCHK, CN_nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_SN_SDFCHK, nCN_D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_SN_SDFCHK, nCN_D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_SN_SDFCHK, nCN_D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_SN_SDFCHK, nCN_nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_SN_SDFCHK, nCN_nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_SN_SDFCHK, nCN_nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSE_SI_SN_SDFCHK, D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SN_SDFCHK, D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nSE_SI_SN_SDFCHK, CN_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nSE_nSI_SN_SDFCHK, CN_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SI_SN_SDFCHK, CN_nD_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SI_SN_SDFCHK, nCN_D_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SI_SN_SDFCHK, nCN_nD_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSI_SN_SDFCHK, CN_D_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSI_nSN_SDFCHK, CN_D_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSI_nSN_SDFCHK, CN_nD_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_D_SE_SN_SDFCHK, CN_D_SE_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSN_SDFCHK, CN_D_SE_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SN_SDFCHK, CN_nD_SE_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSN_SDFCHK, CN_nD_SE_nSN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SN_SDFCHK, nCN_D_SE_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SN_SDFCHK, nCN_nD_SE_SN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    not (nSN, SN);
    and (CN_D_SE_SI_SN, CN, D, SE, SI, SN);
    and (CN_D_SE_SI_nSN, CN, D, SE, SI, nSN);
    and (CN_D_nSE_SI_SN, CN, D, nSE, SI, SN);
    and (CN_D_nSE_SI_nSN, CN, D, nSE, SI, nSN);
    and (CN_D_nSE_nSI_SN, CN, D, nSE, nSI, SN);
    and (CN_D_nSE_nSI_nSN, CN, D, nSE, nSI, nSN);
    and (CN_nD_SE_SI_SN, CN, nD, SE, SI, SN);
    and (CN_nD_SE_SI_nSN, CN, nD, SE, SI, nSN);
    and (CN_nD_nSE_SI_nSN, CN, nD, nSE, SI, nSN);
    and (CN_nD_nSE_nSI_nSN, CN, nD, nSE, nSI, nSN);
    and (nCN_D_SE_SI_SN, nCN, D, SE, SI, SN);
    and (nCN_nD_SE_SI_SN, nCN, nD, SE, SI, SN);
    and (CN_D_SE_nSI_SN, CN, D, SE, nSI, SN);
    and (CN_D_SE_nSI_nSN, CN, D, SE, nSI, nSN);
    and (CN_nD_SE_nSI_SN, CN, nD, SE, nSI, SN);
    and (CN_nD_SE_nSI_nSN, CN, nD, SE, nSI, nSN);
    and (CN_nD_nSE_SI_SN, CN, nD, nSE, SI, SN);
    and (CN_nD_nSE_nSI_SN, CN, nD, nSE, nSI, SN);
    and (nCN_D_SE_nSI_SN, nCN, D, SE, nSI, SN);
    and (nCN_D_nSE_SI_SN, nCN, D, nSE, SI, SN);
    and (nCN_D_nSE_nSI_SN, nCN, D, nSE, nSI, SN);
    and (nCN_nD_SE_nSI_SN, nCN, nD, SE, nSI, SN);
    and (nCN_nD_nSE_SI_SN, nCN, nD, nSE, SI, SN);
    and (nCN_nD_nSE_nSI_SN, nCN, nD, nSE, nSI, SN);
    and (D_nSE_SI_SN, D, nSE, SI, SN);
    and (D_nSE_nSI_SN, D, nSE, nSI, SN);
    and (CN_nSE_SI_SN, CN, nSE, SI, SN);
    and (CN_nSE_nSI_SN, CN, nSE, nSI, SN);
    and (CN_nD_SI_SN, CN, nD, SI, SN);
    and (nCN_D_SI_SN, nCN, D, SI, SN);
    and (nCN_nD_SI_SN, nCN, nD, SI, SN);
    and (CN_D_nSI_SN, CN, D, nSI, SN);
    and (CN_D_nSI_nSN, CN, D, nSI, nSN);
    and (CN_nD_nSI_nSN, CN, nD, nSI, nSN);
    and (CN_D_SE_SN, CN, D, SE, SN);
    and (CN_D_SE_nSN, CN, D, SE, nSN);
    and (CN_nD_SE_SN, CN, nD, SE, SN);
    and (CN_nD_SE_nSN, CN, nD, SE, nSN);
    and (nCN_D_SE_SN, nCN, D, SE, SN);
    and (nCN_nD_SE_SN, nCN, nD, SE, SN);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, CN_d, SN_d);
    and  (SN_check, SE_int_not, CN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, CN, SN);
    and  (SN_check, SE_int_not, CN);
  `endif
  buf  (CN_check, SE_int_not);
   `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& CN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCSNQD0 (SI, D, SE, CP, CN, SN, Q);
    input SI, D, SE, CP, CN, SN;
    output Q;
    reg notifier;
    reg flag;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (DS, S, D_d);
        and (D1, DS, CN_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (DS, S, D);
        and (D1, DS, CN);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 
    buf (CN_i, CN);
    buf (SN_i, SN);
    always @(CN_i or SN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CN_i===1'b0)&&(SN_i===1'b0));
            if (flag == 1) begin 
                if (CN_i!==1'b0) begin
                    $display("%m > CN is released at time %.2fns.", $realtime);
                end 
                if (SN_i!==1'b0) begin
                    $display("%m > SN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CN and SN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SE_SI_SN_SDFCHK, CN_D_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_SI_nSN_SDFCHK, CN_D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SN_SDFCHK, CN_D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_nSN_SDFCHK, CN_D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SN_SDFCHK, CN_D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_nSN_SDFCHK, CN_D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_SN_SDFCHK, CN_nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_nSN_SDFCHK, CN_nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_nSN_SDFCHK, CN_nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_nSN_SDFCHK, CN_nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_SN_SDFCHK, nCN_D_SE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_SN_SDFCHK, nCN_nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_SN_SDFCHK, CN_D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_nSN_SDFCHK, CN_D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_SN_SDFCHK, CN_nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_nSN_SDFCHK, CN_nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SN_SDFCHK, CN_nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SN_SDFCHK, CN_nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_SN_SDFCHK, nCN_D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_SN_SDFCHK, nCN_D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_SN_SDFCHK, nCN_D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_SN_SDFCHK, nCN_nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_SN_SDFCHK, nCN_nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_SN_SDFCHK, nCN_nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSE_SI_SN_SDFCHK, D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SN_SDFCHK, D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nSE_SI_SN_SDFCHK, CN_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nSE_nSI_SN_SDFCHK, CN_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SI_SN_SDFCHK, CN_nD_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SI_SN_SDFCHK, nCN_D_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SI_SN_SDFCHK, nCN_nD_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSI_SN_SDFCHK, CN_D_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSI_nSN_SDFCHK, CN_D_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSI_nSN_SDFCHK, CN_nD_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_D_SE_SN_SDFCHK, CN_D_SE_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSN_SDFCHK, CN_D_SE_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSN_SDFCHK, CN_nD_SE_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SN_SDFCHK, CN_nD_SE_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SN_SDFCHK, nCN_D_SE_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SN_SDFCHK, nCN_nD_SE_SN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    not (nSN, SN);
    and (CN_D_SE_SI_SN, CN, D, SE, SI, SN);
    and (CN_D_SE_SI_nSN, CN, D, SE, SI, nSN);
    and (CN_D_nSE_SI_SN, CN, D, nSE, SI, SN);
    and (CN_D_nSE_SI_nSN, CN, D, nSE, SI, nSN);
    and (CN_D_nSE_nSI_SN, CN, D, nSE, nSI, SN);
    and (CN_D_nSE_nSI_nSN, CN, D, nSE, nSI, nSN);
    and (CN_nD_SE_SI_SN, CN, nD, SE, SI, SN);
    and (CN_nD_SE_SI_nSN, CN, nD, SE, SI, nSN);
    and (CN_nD_nSE_SI_nSN, CN, nD, nSE, SI, nSN);
    and (CN_nD_nSE_nSI_nSN, CN, nD, nSE, nSI, nSN);
    and (nCN_D_SE_SI_SN, nCN, D, SE, SI, SN);
    and (nCN_nD_SE_SI_SN, nCN, nD, SE, SI, SN);
    and (CN_D_SE_nSI_SN, CN, D, SE, nSI, SN);
    and (CN_D_SE_nSI_nSN, CN, D, SE, nSI, nSN);
    and (CN_nD_SE_nSI_SN, CN, nD, SE, nSI, SN);
    and (CN_nD_SE_nSI_nSN, CN, nD, SE, nSI, nSN);
    and (CN_nD_nSE_SI_SN, CN, nD, nSE, SI, SN);
    and (CN_nD_nSE_nSI_SN, CN, nD, nSE, nSI, SN);
    and (nCN_D_SE_nSI_SN, nCN, D, SE, nSI, SN);
    and (nCN_D_nSE_SI_SN, nCN, D, nSE, SI, SN);
    and (nCN_D_nSE_nSI_SN, nCN, D, nSE, nSI, SN);
    and (nCN_nD_SE_nSI_SN, nCN, nD, SE, nSI, SN);
    and (nCN_nD_nSE_SI_SN, nCN, nD, nSE, SI, SN);
    and (nCN_nD_nSE_nSI_SN, nCN, nD, nSE, nSI, SN);
    and (D_nSE_SI_SN, D, nSE, SI, SN);
    and (D_nSE_nSI_SN, D, nSE, nSI, SN);
    and (CN_nSE_SI_SN, CN, nSE, SI, SN);
    and (CN_nSE_nSI_SN, CN, nSE, nSI, SN);
    and (CN_nD_SI_SN, CN, nD, SI, SN);
    and (nCN_D_SI_SN, nCN, D, SI, SN);
    and (nCN_nD_SI_SN, nCN, nD, SI, SN);
    and (CN_D_nSI_SN, CN, D, nSI, SN);
    and (CN_D_nSI_nSN, CN, D, nSI, nSN);
    and (CN_nD_nSI_nSN, CN, nD, nSI, nSN);
    and (CN_D_SE_SN, CN, D, SE, SN);
    and (CN_D_SE_nSN, CN, D, SE, nSN);
    and (CN_nD_SE_nSN, CN, nD, SE, nSN);
    and (CN_nD_SE_SN, CN, nD, SE, SN);
    and (nCN_D_SE_SN, nCN, D, SE, SN);
    and (nCN_nD_SE_SN, nCN, nD, SE, SN);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, CN_d, SN_d);
    and  (SN_check, SE_int_not, CN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, CN, SN);
    and  (SN_check, SE_int_not, CN);
  `endif
  buf  (CN_check, SE_int_not);
   `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& CN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCSNQD1 (SI, D, SE, CP, CN, SN, Q);
    input SI, D, SE, CP, CN, SN;
    output Q;
    reg notifier;
    reg flag;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (DS, S, D_d);
        and (D1, DS, CN_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (DS, S, D);
        and (D1, DS, CN);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 
    buf (CN_i, CN);
    buf (SN_i, SN);
    always @(CN_i or SN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CN_i===1'b0)&&(SN_i===1'b0));
            if (flag == 1) begin 
                if (CN_i!==1'b0) begin
                    $display("%m > CN is released at time %.2fns.", $realtime);
                end 
                if (SN_i!==1'b0) begin
                    $display("%m > SN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CN and SN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SE_SI_SN_SDFCHK, CN_D_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_SI_nSN_SDFCHK, CN_D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SN_SDFCHK, CN_D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_nSN_SDFCHK, CN_D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SN_SDFCHK, CN_D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_nSN_SDFCHK, CN_D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_SN_SDFCHK, CN_nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_nSN_SDFCHK, CN_nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_nSN_SDFCHK, CN_nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_nSN_SDFCHK, CN_nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_SN_SDFCHK, nCN_D_SE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_SN_SDFCHK, nCN_nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_SN_SDFCHK, CN_D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_nSN_SDFCHK, CN_D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_SN_SDFCHK, CN_nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_nSN_SDFCHK, CN_nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SN_SDFCHK, CN_nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SN_SDFCHK, CN_nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_SN_SDFCHK, nCN_D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_SN_SDFCHK, nCN_D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_SN_SDFCHK, nCN_D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_SN_SDFCHK, nCN_nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_SN_SDFCHK, nCN_nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_SN_SDFCHK, nCN_nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSE_SI_SN_SDFCHK, D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SN_SDFCHK, D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nSE_SI_SN_SDFCHK, CN_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nSE_nSI_SN_SDFCHK, CN_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SI_SN_SDFCHK, CN_nD_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SI_SN_SDFCHK, nCN_D_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SI_SN_SDFCHK, nCN_nD_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSI_SN_SDFCHK, CN_D_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSI_nSN_SDFCHK, CN_D_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSI_nSN_SDFCHK, CN_nD_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_D_SE_SN_SDFCHK, CN_D_SE_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSN_SDFCHK, CN_D_SE_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SN_SDFCHK, CN_nD_SE_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSN_SDFCHK, CN_nD_SE_nSN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SN_SDFCHK, nCN_D_SE_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SN_SDFCHK, nCN_nD_SE_SN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    not (nSN, SN);
    and (CN_D_SE_SI_SN, CN, D, SE, SI, SN);
    and (CN_D_SE_SI_nSN, CN, D, SE, SI, nSN);
    and (CN_D_nSE_SI_SN, CN, D, nSE, SI, SN);
    and (CN_D_nSE_SI_nSN, CN, D, nSE, SI, nSN);
    and (CN_D_nSE_nSI_SN, CN, D, nSE, nSI, SN);
    and (CN_D_nSE_nSI_nSN, CN, D, nSE, nSI, nSN);
    and (CN_nD_SE_SI_SN, CN, nD, SE, SI, SN);
    and (CN_nD_SE_SI_nSN, CN, nD, SE, SI, nSN);
    and (CN_nD_nSE_SI_nSN, CN, nD, nSE, SI, nSN);
    and (CN_nD_nSE_nSI_nSN, CN, nD, nSE, nSI, nSN);
    and (nCN_D_SE_SI_SN, nCN, D, SE, SI, SN);
    and (nCN_nD_SE_SI_SN, nCN, nD, SE, SI, SN);
    and (CN_D_SE_nSI_SN, CN, D, SE, nSI, SN);
    and (CN_D_SE_nSI_nSN, CN, D, SE, nSI, nSN);
    and (CN_nD_SE_nSI_SN, CN, nD, SE, nSI, SN);
    and (CN_nD_SE_nSI_nSN, CN, nD, SE, nSI, nSN);
    and (CN_nD_nSE_SI_SN, CN, nD, nSE, SI, SN);
    and (CN_nD_nSE_nSI_SN, CN, nD, nSE, nSI, SN);
    and (nCN_D_SE_nSI_SN, nCN, D, SE, nSI, SN);
    and (nCN_D_nSE_SI_SN, nCN, D, nSE, SI, SN);
    and (nCN_D_nSE_nSI_SN, nCN, D, nSE, nSI, SN);
    and (nCN_nD_SE_nSI_SN, nCN, nD, SE, nSI, SN);
    and (nCN_nD_nSE_SI_SN, nCN, nD, nSE, SI, SN);
    and (nCN_nD_nSE_nSI_SN, nCN, nD, nSE, nSI, SN);
    and (D_nSE_SI_SN, D, nSE, SI, SN);
    and (D_nSE_nSI_SN, D, nSE, nSI, SN);
    and (CN_nSE_SI_SN, CN, nSE, SI, SN);
    and (CN_nSE_nSI_SN, CN, nSE, nSI, SN);
    and (CN_nD_SI_SN, CN, nD, SI, SN);
    and (nCN_D_SI_SN, nCN, D, SI, SN);
    and (nCN_nD_SI_SN, nCN, nD, SI, SN);
    and (CN_D_nSI_SN, CN, D, nSI, SN);
    and (CN_D_nSI_nSN, CN, D, nSI, nSN);
    and (CN_nD_nSI_nSN, CN, nD, nSI, nSN);
    and (CN_D_SE_SN, CN, D, SE, SN);
    and (CN_D_SE_nSN, CN, D, SE, nSN);
    and (CN_nD_SE_SN, CN, nD, SE, SN);
    and (CN_nD_SE_nSN, CN, nD, SE, nSN);
    and (nCN_D_SE_SN, nCN, D, SE, SN);
    and (nCN_nD_SE_SN, nCN, nD, SE, SN);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, CN_d, SN_d);
    and  (SN_check, SE_int_not, CN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, CN, SN);
    and  (SN_check, SE_int_not, CN);
  `endif
  buf  (CN_check, SE_int_not);
   `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& CN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCSNQD2 (SI, D, SE, CP, CN, SN, Q);
    input SI, D, SE, CP, CN, SN;
    output Q;
    reg notifier;
    reg flag;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (DS, S, D_d);
        and (D1, DS, CN_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (DS, S, D);
        and (D1, DS, CN);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 
    buf (CN_i, CN);
    buf (SN_i, SN);
    always @(CN_i or SN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CN_i===1'b0)&&(SN_i===1'b0));
            if (flag == 1) begin 
                if (CN_i!==1'b0) begin
                    $display("%m > CN is released at time %.2fns.", $realtime);
                end 
                if (SN_i!==1'b0) begin
                    $display("%m > SN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CN and SN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SE_SI_SN_SDFCHK, CN_D_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_SI_nSN_SDFCHK, CN_D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SN_SDFCHK, CN_D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_nSN_SDFCHK, CN_D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SN_SDFCHK, CN_D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_nSN_SDFCHK, CN_D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_SN_SDFCHK, CN_nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_nSN_SDFCHK, CN_nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_nSN_SDFCHK, CN_nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_nSN_SDFCHK, CN_nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_SN_SDFCHK, nCN_D_SE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_SN_SDFCHK, nCN_nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_SN_SDFCHK, CN_D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_nSN_SDFCHK, CN_D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_SN_SDFCHK, CN_nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_nSN_SDFCHK, CN_nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SN_SDFCHK, CN_nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SN_SDFCHK, CN_nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_SN_SDFCHK, nCN_D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_SN_SDFCHK, nCN_D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_SN_SDFCHK, nCN_D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_SN_SDFCHK, nCN_nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_SN_SDFCHK, nCN_nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_SN_SDFCHK, nCN_nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSE_SI_SN_SDFCHK, D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SN_SDFCHK, D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nSE_SI_SN_SDFCHK, CN_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nSE_nSI_SN_SDFCHK, CN_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SI_SN_SDFCHK, CN_nD_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SI_SN_SDFCHK, nCN_D_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SI_SN_SDFCHK, nCN_nD_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSI_SN_SDFCHK, CN_D_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSI_nSN_SDFCHK, CN_D_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSI_nSN_SDFCHK, CN_nD_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_D_SE_SN_SDFCHK, CN_D_SE_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSN_SDFCHK, CN_D_SE_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SN_SDFCHK, CN_nD_SE_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSN_SDFCHK, CN_nD_SE_nSN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SN_SDFCHK, nCN_D_SE_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SN_SDFCHK, nCN_nD_SE_SN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    not (nSN, SN);
    and (CN_D_SE_SI_SN, CN, D, SE, SI, SN);
    and (CN_D_SE_SI_nSN, CN, D, SE, SI, nSN);
    and (CN_D_nSE_SI_SN, CN, D, nSE, SI, SN);
    and (CN_D_nSE_SI_nSN, CN, D, nSE, SI, nSN);
    and (CN_D_nSE_nSI_SN, CN, D, nSE, nSI, SN);
    and (CN_D_nSE_nSI_nSN, CN, D, nSE, nSI, nSN);
    and (CN_nD_SE_SI_SN, CN, nD, SE, SI, SN);
    and (CN_nD_SE_SI_nSN, CN, nD, SE, SI, nSN);
    and (CN_nD_nSE_SI_nSN, CN, nD, nSE, SI, nSN);
    and (CN_nD_nSE_nSI_nSN, CN, nD, nSE, nSI, nSN);
    and (nCN_D_SE_SI_SN, nCN, D, SE, SI, SN);
    and (nCN_nD_SE_SI_SN, nCN, nD, SE, SI, SN);
    and (CN_D_SE_nSI_SN, CN, D, SE, nSI, SN);
    and (CN_D_SE_nSI_nSN, CN, D, SE, nSI, nSN);
    and (CN_nD_SE_nSI_SN, CN, nD, SE, nSI, SN);
    and (CN_nD_SE_nSI_nSN, CN, nD, SE, nSI, nSN);
    and (CN_nD_nSE_SI_SN, CN, nD, nSE, SI, SN);
    and (CN_nD_nSE_nSI_SN, CN, nD, nSE, nSI, SN);
    and (nCN_D_SE_nSI_SN, nCN, D, SE, nSI, SN);
    and (nCN_D_nSE_SI_SN, nCN, D, nSE, SI, SN);
    and (nCN_D_nSE_nSI_SN, nCN, D, nSE, nSI, SN);
    and (nCN_nD_SE_nSI_SN, nCN, nD, SE, nSI, SN);
    and (nCN_nD_nSE_SI_SN, nCN, nD, nSE, SI, SN);
    and (nCN_nD_nSE_nSI_SN, nCN, nD, nSE, nSI, SN);
    and (D_nSE_SI_SN, D, nSE, SI, SN);
    and (D_nSE_nSI_SN, D, nSE, nSI, SN);
    and (CN_nSE_SI_SN, CN, nSE, SI, SN);
    and (CN_nSE_nSI_SN, CN, nSE, nSI, SN);
    and (CN_nD_SI_SN, CN, nD, SI, SN);
    and (nCN_D_SI_SN, nCN, D, SI, SN);
    and (nCN_nD_SI_SN, nCN, nD, SI, SN);
    and (CN_D_nSI_SN, CN, D, nSI, SN);
    and (CN_D_nSI_nSN, CN, D, nSI, nSN);
    and (CN_nD_nSI_nSN, CN, nD, nSI, nSN);
    and (CN_D_SE_SN, CN, D, SE, SN);
    and (CN_D_SE_nSN, CN, D, SE, nSN);
    and (CN_nD_SE_SN, CN, nD, SE, SN);
    and (CN_nD_SE_nSN, CN, nD, SE, nSN);
    and (nCN_D_SE_SN, nCN, D, SE, SN);
    and (nCN_nD_SE_SN, nCN, nD, SE, SN);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, CN_d, SN_d);
    and  (SN_check, SE_int_not, CN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, CN, SN);
    and  (SN_check, SE_int_not, CN);
  `endif
  buf  (CN_check, SE_int_not);
   `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& CN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCSNQD4 (SI, D, SE, CP, CN, SN, Q);
    input SI, D, SE, CP, CN, SN;
    output Q;
    reg notifier;
    reg flag;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (DS, S, D_d);
        and (D1, DS, CN_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (DS, S, D);
        and (D1, DS, CN);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 
    buf (CN_i, CN);
    buf (SN_i, SN);
    always @(CN_i or SN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CN_i===1'b0)&&(SN_i===1'b0));
            if (flag == 1) begin 
                if (CN_i!==1'b0) begin
                    $display("%m > CN is released at time %.2fns.", $realtime);
                end 
                if (SN_i!==1'b0) begin
                    $display("%m > SN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CN and SN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SE_SI_SN_SDFCHK, CN_D_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_SI_nSN_SDFCHK, CN_D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SN_SDFCHK, CN_D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_nSN_SDFCHK, CN_D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SN_SDFCHK, CN_D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_nSN_SDFCHK, CN_D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_SN_SDFCHK, CN_nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_nSN_SDFCHK, CN_nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_nSN_SDFCHK, CN_nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_nSN_SDFCHK, CN_nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_SN_SDFCHK, nCN_D_SE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_SN_SDFCHK, nCN_nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_SN_SDFCHK, CN_D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_nSN_SDFCHK, CN_D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_SN_SDFCHK, CN_nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_nSN_SDFCHK, CN_nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SN_SDFCHK, CN_nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SN_SDFCHK, CN_nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_SN_SDFCHK, nCN_D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_SN_SDFCHK, nCN_D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_SN_SDFCHK, nCN_D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_SN_SDFCHK, nCN_nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_SN_SDFCHK, nCN_nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_SN_SDFCHK, nCN_nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSE_SI_SN_SDFCHK, D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SN_SDFCHK, D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nSE_SI_SN_SDFCHK, CN_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nSE_nSI_SN_SDFCHK, CN_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SI_SN_SDFCHK, CN_nD_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SI_SN_SDFCHK, nCN_D_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SI_SN_SDFCHK, nCN_nD_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSI_SN_SDFCHK, CN_D_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSI_nSN_SDFCHK, CN_D_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSI_nSN_SDFCHK, CN_nD_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_D_SE_SN_SDFCHK, CN_D_SE_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSN_SDFCHK, CN_D_SE_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SN_SDFCHK, CN_nD_SE_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSN_SDFCHK, CN_nD_SE_nSN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SN_SDFCHK, nCN_D_SE_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SN_SDFCHK, nCN_nD_SE_SN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    not (nSN, SN);
    and (CN_D_SE_SI_SN, CN, D, SE, SI, SN);
    and (CN_D_SE_SI_nSN, CN, D, SE, SI, nSN);
    and (CN_D_nSE_SI_SN, CN, D, nSE, SI, SN);
    and (CN_D_nSE_SI_nSN, CN, D, nSE, SI, nSN);
    and (CN_D_nSE_nSI_SN, CN, D, nSE, nSI, SN);
    and (CN_D_nSE_nSI_nSN, CN, D, nSE, nSI, nSN);
    and (CN_nD_SE_SI_SN, CN, nD, SE, SI, SN);
    and (CN_nD_SE_SI_nSN, CN, nD, SE, SI, nSN);
    and (CN_nD_nSE_SI_nSN, CN, nD, nSE, SI, nSN);
    and (CN_nD_nSE_nSI_nSN, CN, nD, nSE, nSI, nSN);
    and (nCN_D_SE_SI_SN, nCN, D, SE, SI, SN);
    and (nCN_nD_SE_SI_SN, nCN, nD, SE, SI, SN);
    and (CN_D_SE_nSI_SN, CN, D, SE, nSI, SN);
    and (CN_D_SE_nSI_nSN, CN, D, SE, nSI, nSN);
    and (CN_nD_SE_nSI_SN, CN, nD, SE, nSI, SN);
    and (CN_nD_SE_nSI_nSN, CN, nD, SE, nSI, nSN);
    and (CN_nD_nSE_SI_SN, CN, nD, nSE, SI, SN);
    and (CN_nD_nSE_nSI_SN, CN, nD, nSE, nSI, SN);
    and (nCN_D_SE_nSI_SN, nCN, D, SE, nSI, SN);
    and (nCN_D_nSE_SI_SN, nCN, D, nSE, SI, SN);
    and (nCN_D_nSE_nSI_SN, nCN, D, nSE, nSI, SN);
    and (nCN_nD_SE_nSI_SN, nCN, nD, SE, nSI, SN);
    and (nCN_nD_nSE_SI_SN, nCN, nD, nSE, SI, SN);
    and (nCN_nD_nSE_nSI_SN, nCN, nD, nSE, nSI, SN);
    and (D_nSE_SI_SN, D, nSE, SI, SN);
    and (D_nSE_nSI_SN, D, nSE, nSI, SN);
    and (CN_nSE_SI_SN, CN, nSE, SI, SN);
    and (CN_nSE_nSI_SN, CN, nSE, nSI, SN);
    and (CN_nD_SI_SN, CN, nD, SI, SN);
    and (nCN_D_SI_SN, nCN, D, SI, SN);
    and (nCN_nD_SI_SN, nCN, nD, SI, SN);
    and (CN_D_nSI_SN, CN, D, nSI, SN);
    and (CN_D_nSI_nSN, CN, D, nSI, nSN);
    and (CN_nD_nSI_nSN, CN, nD, nSI, nSN);
    and (CN_D_SE_SN, CN, D, SE, SN);
    and (CN_D_SE_nSN, CN, D, SE, nSN);
    and (CN_nD_SE_SN, CN, nD, SE, SN);
    and (CN_nD_SE_nSN, CN, nD, SE, nSN);
    and (nCN_D_SE_SN, nCN, D, SE, SN);
    and (nCN_nD_SE_SN, nCN, nD, SE, SN);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, CN_d, SN_d);
    and  (SN_check, SE_int_not, CN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, CN, SN);
    and  (SN_check, SE_int_not, CN);
  `endif
  buf  (CN_check, SE_int_not);
   `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& CN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKSND0 (SI, D, SE, CP, SN, Q, QN);
    input SI, D, SE, CP, SN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (D1, S, D_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (D1, S, D);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SN_SDFCHK, D_SE_SI_SN, 1'b1);
    tsmc_xbuf (D_SE_SI_nSN_SDFCHK, D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_SI_SN_SDFCHK, D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (D_nSE_SI_nSN_SDFCHK, D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SN_SDFCHK, D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_nSN_SDFCHK, D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_SE_SI_SN_SDFCHK, nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (nD_SE_SI_nSN_SDFCHK, nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_nSN_SDFCHK, nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_nSN_SDFCHK, nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (D_SE_nSI_SN_SDFCHK, D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (D_SE_nSI_nSN_SDFCHK, D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SN_SDFCHK, nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nD_SE_nSI_nSN_SDFCHK, nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SN_SDFCHK, nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SN_SDFCHK, nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nSE_SI_SN_SDFCHK, nSE_SI_SN, 1'b1);
    tsmc_xbuf (nSE_nSI_SN_SDFCHK, nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nD_SI_SN_SDFCHK, nD_SI_SN, 1'b1);
    tsmc_xbuf (D_nSI_SN_SDFCHK, D_nSI_SN, 1'b1);
    tsmc_xbuf (nD_nSI_nSN_SDFCHK, nD_nSI_nSN, 1'b1);
    tsmc_xbuf (D_nSI_nSN_SDFCHK, D_nSI_nSN, 1'b1);
    tsmc_xbuf (D_SE_SN_SDFCHK, D_SE_SN, 1'b1);
    tsmc_xbuf (D_SE_nSN_SDFCHK, D_SE_nSN, 1'b1);
    tsmc_xbuf (nD_SE_SN_SDFCHK, nD_SE_SN, 1'b1);
    tsmc_xbuf (nD_SE_nSN_SDFCHK, nD_SE_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nSN, SN);
    and (D_SE_SI_SN, D, SE, SI, SN);
    and (D_SE_SI_nSN, D, SE, SI, nSN);
    and (D_nSE_SI_SN, D, nSE, SI, SN);
    and (D_nSE_SI_nSN, D, nSE, SI, nSN);
    and (D_nSE_nSI_SN, D, nSE, nSI, SN);
    and (D_nSE_nSI_nSN, D, nSE, nSI, nSN);
    and (nD_SE_SI_SN, nD, SE, SI, SN);
    and (nD_SE_SI_nSN, nD, SE, SI, nSN);
    and (nD_nSE_SI_nSN, nD, nSE, SI, nSN);
    and (nD_nSE_nSI_nSN, nD, nSE, nSI, nSN);
    and (D_SE_nSI_SN, D, SE, nSI, SN);
    and (D_SE_nSI_nSN, D, SE, nSI, nSN);
    and (nD_SE_nSI_SN, nD, SE, nSI, SN);
    and (nD_SE_nSI_nSN, nD, SE, nSI, nSN);
    and (nD_nSE_SI_SN, nD, nSE, SI, SN);
    and (nD_nSE_nSI_SN, nD, nSE, nSI, SN);
    and (nSE_SI_SN, nSE, SI, SN);
    and (nSE_nSI_SN, nSE, nSI, SN);
    and (nD_SI_SN, nD, SI, SN);
    and (D_nSI_SN, D, nSI, SN);
    and (nD_nSI_nSN, nD, nSI, nSN);
    and (D_nSI_nSN, D, nSI, nSN);
    and (D_SE_SN, D, SE, SN);
    and (D_SE_nSN, D, SE, nSN);
    and (nD_SE_SN, nD, SE, SN);
    and (nD_SE_nSN, nD, SE, nSN);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, SN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, SN);
  `endif
  buf  (SN_check, SE_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKSND1 (SI, D, SE, CP, SN, Q, QN);
    input SI, D, SE, CP, SN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (D1, S, D_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (D1, S, D);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SN_SDFCHK, D_SE_SI_SN, 1'b1);
    tsmc_xbuf (D_SE_SI_nSN_SDFCHK, D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_SI_SN_SDFCHK, D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (D_nSE_SI_nSN_SDFCHK, D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SN_SDFCHK, D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_nSN_SDFCHK, D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_SE_SI_SN_SDFCHK, nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (nD_SE_SI_nSN_SDFCHK, nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_nSN_SDFCHK, nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_nSN_SDFCHK, nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (D_SE_nSI_SN_SDFCHK, D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (D_SE_nSI_nSN_SDFCHK, D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SN_SDFCHK, nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nD_SE_nSI_nSN_SDFCHK, nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SN_SDFCHK, nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SN_SDFCHK, nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nSE_SI_SN_SDFCHK, nSE_SI_SN, 1'b1);
    tsmc_xbuf (nSE_nSI_SN_SDFCHK, nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nD_SI_SN_SDFCHK, nD_SI_SN, 1'b1);
    tsmc_xbuf (D_nSI_SN_SDFCHK, D_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSI_nSN_SDFCHK, D_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_nSI_nSN_SDFCHK, nD_nSI_nSN, 1'b1);
    tsmc_xbuf (D_SE_SN_SDFCHK, D_SE_SN, 1'b1);
    tsmc_xbuf (D_SE_nSN_SDFCHK, D_SE_nSN, 1'b1);
    tsmc_xbuf (nD_SE_SN_SDFCHK, nD_SE_SN, 1'b1);
    tsmc_xbuf (nD_SE_nSN_SDFCHK, nD_SE_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nSN, SN);
    and (D_SE_SI_SN, D, SE, SI, SN);
    and (D_SE_SI_nSN, D, SE, SI, nSN);
    and (D_nSE_SI_SN, D, nSE, SI, SN);
    and (D_nSE_SI_nSN, D, nSE, SI, nSN);
    and (D_nSE_nSI_SN, D, nSE, nSI, SN);
    and (D_nSE_nSI_nSN, D, nSE, nSI, nSN);
    and (nD_SE_SI_SN, nD, SE, SI, SN);
    and (nD_SE_SI_nSN, nD, SE, SI, nSN);
    and (nD_nSE_SI_nSN, nD, nSE, SI, nSN);
    and (nD_nSE_nSI_nSN, nD, nSE, nSI, nSN);
    and (D_SE_nSI_SN, D, SE, nSI, SN);
    and (D_SE_nSI_nSN, D, SE, nSI, nSN);
    and (nD_SE_nSI_SN, nD, SE, nSI, SN);
    and (nD_SE_nSI_nSN, nD, SE, nSI, nSN);
    and (nD_nSE_SI_SN, nD, nSE, SI, SN);
    and (nD_nSE_nSI_SN, nD, nSE, nSI, SN);
    and (nSE_SI_SN, nSE, SI, SN);
    and (nSE_nSI_SN, nSE, nSI, SN);
    and (nD_SI_SN, nD, SI, SN);
    and (D_nSI_SN, D, nSI, SN);
    and (D_nSI_nSN, D, nSI, nSN);
    and (nD_nSI_nSN, nD, nSI, nSN);
    and (D_SE_SN, D, SE, SN);
    and (D_SE_nSN, D, SE, nSN);
    and (nD_SE_SN, nD, SE, SN);
    and (nD_SE_nSN, nD, SE, nSN);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, SN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, SN);
  `endif
  buf  (SN_check, SE_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKSND2 (SI, D, SE, CP, SN, Q, QN);
    input SI, D, SE, CP, SN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (D1, S, D_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (D1, S, D);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SN_SDFCHK, D_SE_SI_SN, 1'b1);
    tsmc_xbuf (D_SE_SI_nSN_SDFCHK, D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_SI_SN_SDFCHK, D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (D_nSE_SI_nSN_SDFCHK, D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SN_SDFCHK, D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_nSN_SDFCHK, D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_SE_SI_SN_SDFCHK, nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (nD_SE_SI_nSN_SDFCHK, nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_nSN_SDFCHK, nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_nSN_SDFCHK, nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (D_SE_nSI_SN_SDFCHK, D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (D_SE_nSI_nSN_SDFCHK, D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SN_SDFCHK, nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nD_SE_nSI_nSN_SDFCHK, nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SN_SDFCHK, nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SN_SDFCHK, nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nSE_SI_SN_SDFCHK, nSE_SI_SN, 1'b1);
    tsmc_xbuf (nSE_nSI_SN_SDFCHK, nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nD_SI_SN_SDFCHK, nD_SI_SN, 1'b1);
    tsmc_xbuf (D_nSI_SN_SDFCHK, D_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSI_nSN_SDFCHK, D_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_nSI_nSN_SDFCHK, nD_nSI_nSN, 1'b1);
    tsmc_xbuf (D_SE_SN_SDFCHK, D_SE_SN, 1'b1);
    tsmc_xbuf (D_SE_nSN_SDFCHK, D_SE_nSN, 1'b1);
    tsmc_xbuf (nD_SE_SN_SDFCHK, nD_SE_SN, 1'b1);
    tsmc_xbuf (nD_SE_nSN_SDFCHK, nD_SE_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nSN, SN);
    and (D_SE_SI_SN, D, SE, SI, SN);
    and (D_SE_SI_nSN, D, SE, SI, nSN);
    and (D_nSE_SI_SN, D, nSE, SI, SN);
    and (D_nSE_SI_nSN, D, nSE, SI, nSN);
    and (D_nSE_nSI_SN, D, nSE, nSI, SN);
    and (D_nSE_nSI_nSN, D, nSE, nSI, nSN);
    and (nD_SE_SI_SN, nD, SE, SI, SN);
    and (nD_SE_SI_nSN, nD, SE, SI, nSN);
    and (nD_nSE_SI_nSN, nD, nSE, SI, nSN);
    and (nD_nSE_nSI_nSN, nD, nSE, nSI, nSN);
    and (D_SE_nSI_SN, D, SE, nSI, SN);
    and (D_SE_nSI_nSN, D, SE, nSI, nSN);
    and (nD_SE_nSI_SN, nD, SE, nSI, SN);
    and (nD_SE_nSI_nSN, nD, SE, nSI, nSN);
    and (nD_nSE_SI_SN, nD, nSE, SI, SN);
    and (nD_nSE_nSI_SN, nD, nSE, nSI, SN);
    and (nSE_SI_SN, nSE, SI, SN);
    and (nSE_nSI_SN, nSE, nSI, SN);
    and (nD_SI_SN, nD, SI, SN);
    and (D_nSI_SN, D, nSI, SN);
    and (D_nSI_nSN, D, nSI, nSN);
    and (nD_nSI_nSN, nD, nSI, nSN);
    and (D_SE_SN, D, SE, SN);
    and (D_SE_nSN, D, SE, nSN);
    and (nD_SE_SN, nD, SE, SN);
    and (nD_SE_nSN, nD, SE, nSN);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, SN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, SN);
  `endif
  buf  (SN_check, SE_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKSND4 (SI, D, SE, CP, SN, Q, QN);
    input SI, D, SE, CP, SN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (D1, S, D_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (D1, S, D);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SN_SDFCHK, D_SE_SI_SN, 1'b1);
    tsmc_xbuf (D_SE_SI_nSN_SDFCHK, D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_SI_SN_SDFCHK, D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (D_nSE_SI_nSN_SDFCHK, D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SN_SDFCHK, D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_nSN_SDFCHK, D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_SE_SI_SN_SDFCHK, nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (nD_SE_SI_nSN_SDFCHK, nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_nSN_SDFCHK, nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_nSN_SDFCHK, nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (D_SE_nSI_SN_SDFCHK, D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (D_SE_nSI_nSN_SDFCHK, D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SN_SDFCHK, nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nD_SE_nSI_nSN_SDFCHK, nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SN_SDFCHK, nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SN_SDFCHK, nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nSE_SI_SN_SDFCHK, nSE_SI_SN, 1'b1);
    tsmc_xbuf (nSE_nSI_SN_SDFCHK, nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nD_SI_SN_SDFCHK, nD_SI_SN, 1'b1);
    tsmc_xbuf (D_nSI_SN_SDFCHK, D_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSI_nSN_SDFCHK, D_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_nSI_nSN_SDFCHK, nD_nSI_nSN, 1'b1);
    tsmc_xbuf (D_SE_SN_SDFCHK, D_SE_SN, 1'b1);
    tsmc_xbuf (D_SE_nSN_SDFCHK, D_SE_nSN, 1'b1);
    tsmc_xbuf (nD_SE_SN_SDFCHK, nD_SE_SN, 1'b1);
    tsmc_xbuf (nD_SE_nSN_SDFCHK, nD_SE_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nSN, SN);
    and (D_SE_SI_SN, D, SE, SI, SN);
    and (D_SE_SI_nSN, D, SE, SI, nSN);
    and (D_nSE_SI_SN, D, nSE, SI, SN);
    and (D_nSE_SI_nSN, D, nSE, SI, nSN);
    and (D_nSE_nSI_SN, D, nSE, nSI, SN);
    and (D_nSE_nSI_nSN, D, nSE, nSI, nSN);
    and (nD_SE_SI_SN, nD, SE, SI, SN);
    and (nD_SE_SI_nSN, nD, SE, SI, nSN);
    and (nD_nSE_SI_nSN, nD, nSE, SI, nSN);
    and (nD_nSE_nSI_nSN, nD, nSE, nSI, nSN);
    and (D_SE_nSI_SN, D, SE, nSI, SN);
    and (D_SE_nSI_nSN, D, SE, nSI, nSN);
    and (nD_SE_nSI_SN, nD, SE, nSI, SN);
    and (nD_SE_nSI_nSN, nD, SE, nSI, nSN);
    and (nD_nSE_SI_SN, nD, nSE, SI, SN);
    and (nD_nSE_nSI_SN, nD, nSE, nSI, SN);
    and (nSE_SI_SN, nSE, SI, SN);
    and (nSE_nSI_SN, nSE, nSI, SN);
    and (nD_SI_SN, nD, SI, SN);
    and (D_nSI_SN, D, nSI, SN);
    and (D_nSI_nSN, D, nSI, nSN);
    and (nD_nSI_nSN, nD, nSI, nSN);
    and (D_SE_SN, D, SE, SN);
    and (D_SE_nSN, D, SE, nSN);
    and (nD_SE_SN, nD, SE, SN);
    and (nD_SE_nSN, nD, SE, nSN);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, SN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, SN);
  `endif
  buf  (SN_check, SE_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKSNQD0 (SI, D, SE, CP, SN, Q);
    input SI, D, SE, CP, SN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (D1, S, D_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (D1, S, D);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SN_SDFCHK, D_SE_SI_SN, 1'b1);
    tsmc_xbuf (D_SE_SI_nSN_SDFCHK, D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_SI_SN_SDFCHK, D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (D_nSE_SI_nSN_SDFCHK, D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SN_SDFCHK, D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_nSN_SDFCHK, D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_SE_SI_SN_SDFCHK, nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (nD_SE_SI_nSN_SDFCHK, nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_nSN_SDFCHK, nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_nSN_SDFCHK, nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (D_SE_nSI_SN_SDFCHK, D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (D_SE_nSI_nSN_SDFCHK, D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SN_SDFCHK, nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nD_SE_nSI_nSN_SDFCHK, nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SN_SDFCHK, nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SN_SDFCHK, nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nSE_SI_SN_SDFCHK, nSE_SI_SN, 1'b1);
    tsmc_xbuf (nSE_nSI_SN_SDFCHK, nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nD_SI_SN_SDFCHK, nD_SI_SN, 1'b1);
    tsmc_xbuf (D_nSI_SN_SDFCHK, D_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSI_nSN_SDFCHK, D_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_nSI_nSN_SDFCHK, nD_nSI_nSN, 1'b1);
    tsmc_xbuf (D_SE_SN_SDFCHK, D_SE_SN, 1'b1);
    tsmc_xbuf (D_SE_nSN_SDFCHK, D_SE_nSN, 1'b1);
    tsmc_xbuf (nD_SE_nSN_SDFCHK, nD_SE_nSN, 1'b1);
    tsmc_xbuf (nD_SE_SN_SDFCHK, nD_SE_SN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nSN, SN);
    and (D_SE_SI_SN, D, SE, SI, SN);
    and (D_SE_SI_nSN, D, SE, SI, nSN);
    and (D_nSE_SI_SN, D, nSE, SI, SN);
    and (D_nSE_SI_nSN, D, nSE, SI, nSN);
    and (D_nSE_nSI_SN, D, nSE, nSI, SN);
    and (D_nSE_nSI_nSN, D, nSE, nSI, nSN);
    and (nD_SE_SI_SN, nD, SE, SI, SN);
    and (nD_SE_SI_nSN, nD, SE, SI, nSN);
    and (nD_nSE_SI_nSN, nD, nSE, SI, nSN);
    and (nD_nSE_nSI_nSN, nD, nSE, nSI, nSN);
    and (D_SE_nSI_SN, D, SE, nSI, SN);
    and (D_SE_nSI_nSN, D, SE, nSI, nSN);
    and (nD_SE_nSI_SN, nD, SE, nSI, SN);
    and (nD_SE_nSI_nSN, nD, SE, nSI, nSN);
    and (nD_nSE_SI_SN, nD, nSE, SI, SN);
    and (nD_nSE_nSI_SN, nD, nSE, nSI, SN);
    and (nSE_SI_SN, nSE, SI, SN);
    and (nSE_nSI_SN, nSE, nSI, SN);
    and (nD_SI_SN, nD, SI, SN);
    and (D_nSI_SN, D, nSI, SN);
    and (D_nSI_nSN, D, nSI, nSN);
    and (nD_nSI_nSN, nD, nSI, nSN);
    and (D_SE_SN, D, SE, SN);
    and (D_SE_nSN, D, SE, nSN);
    and (nD_SE_nSN, nD, SE, nSN);
    and (nD_SE_SN, nD, SE, SN);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, SN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, SN);
  `endif
  buf  (SN_check, SE_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKSNQD1 (SI, D, SE, CP, SN, Q);
    input SI, D, SE, CP, SN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (D1, S, D_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (D1, S, D);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SN_SDFCHK, D_SE_SI_SN, 1'b1);
    tsmc_xbuf (D_SE_SI_nSN_SDFCHK, D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_SI_SN_SDFCHK, D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (D_nSE_SI_nSN_SDFCHK, D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SN_SDFCHK, D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_nSN_SDFCHK, D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_SE_SI_SN_SDFCHK, nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (nD_SE_SI_nSN_SDFCHK, nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_nSN_SDFCHK, nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_nSN_SDFCHK, nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (D_SE_nSI_SN_SDFCHK, D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (D_SE_nSI_nSN_SDFCHK, D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SN_SDFCHK, nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nD_SE_nSI_nSN_SDFCHK, nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SN_SDFCHK, nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SN_SDFCHK, nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nSE_SI_SN_SDFCHK, nSE_SI_SN, 1'b1);
    tsmc_xbuf (nSE_nSI_SN_SDFCHK, nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nD_SI_SN_SDFCHK, nD_SI_SN, 1'b1);
    tsmc_xbuf (D_nSI_SN_SDFCHK, D_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSI_nSN_SDFCHK, D_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_nSI_nSN_SDFCHK, nD_nSI_nSN, 1'b1);
    tsmc_xbuf (D_SE_SN_SDFCHK, D_SE_SN, 1'b1);
    tsmc_xbuf (D_SE_nSN_SDFCHK, D_SE_nSN, 1'b1);
    tsmc_xbuf (nD_SE_SN_SDFCHK, nD_SE_SN, 1'b1);
    tsmc_xbuf (nD_SE_nSN_SDFCHK, nD_SE_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nSN, SN);
    and (D_SE_SI_SN, D, SE, SI, SN);
    and (D_SE_SI_nSN, D, SE, SI, nSN);
    and (D_nSE_SI_SN, D, nSE, SI, SN);
    and (D_nSE_SI_nSN, D, nSE, SI, nSN);
    and (D_nSE_nSI_SN, D, nSE, nSI, SN);
    and (D_nSE_nSI_nSN, D, nSE, nSI, nSN);
    and (nD_SE_SI_SN, nD, SE, SI, SN);
    and (nD_SE_SI_nSN, nD, SE, SI, nSN);
    and (nD_nSE_SI_nSN, nD, nSE, SI, nSN);
    and (nD_nSE_nSI_nSN, nD, nSE, nSI, nSN);
    and (D_SE_nSI_SN, D, SE, nSI, SN);
    and (D_SE_nSI_nSN, D, SE, nSI, nSN);
    and (nD_SE_nSI_SN, nD, SE, nSI, SN);
    and (nD_SE_nSI_nSN, nD, SE, nSI, nSN);
    and (nD_nSE_SI_SN, nD, nSE, SI, SN);
    and (nD_nSE_nSI_SN, nD, nSE, nSI, SN);
    and (nSE_SI_SN, nSE, SI, SN);
    and (nSE_nSI_SN, nSE, nSI, SN);
    and (nD_SI_SN, nD, SI, SN);
    and (D_nSI_SN, D, nSI, SN);
    and (D_nSI_nSN, D, nSI, nSN);
    and (nD_nSI_nSN, nD, nSI, nSN);
    and (D_SE_SN, D, SE, SN);
    and (D_SE_nSN, D, SE, nSN);
    and (nD_SE_SN, nD, SE, SN);
    and (nD_SE_nSN, nD, SE, nSN);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, SN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, SN);
  `endif
  buf  (SN_check, SE_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKSNQD2 (SI, D, SE, CP, SN, Q);
    input SI, D, SE, CP, SN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (D1, S, D_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (D1, S, D);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SN_SDFCHK, D_SE_SI_SN, 1'b1);
    tsmc_xbuf (D_SE_SI_nSN_SDFCHK, D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_SI_SN_SDFCHK, D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (D_nSE_SI_nSN_SDFCHK, D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SN_SDFCHK, D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_nSN_SDFCHK, D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_SE_SI_SN_SDFCHK, nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (nD_SE_SI_nSN_SDFCHK, nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_nSN_SDFCHK, nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_nSN_SDFCHK, nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (D_SE_nSI_SN_SDFCHK, D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (D_SE_nSI_nSN_SDFCHK, D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SN_SDFCHK, nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nD_SE_nSI_nSN_SDFCHK, nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SN_SDFCHK, nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SN_SDFCHK, nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nSE_SI_SN_SDFCHK, nSE_SI_SN, 1'b1);
    tsmc_xbuf (nSE_nSI_SN_SDFCHK, nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nD_SI_SN_SDFCHK, nD_SI_SN, 1'b1);
    tsmc_xbuf (D_nSI_SN_SDFCHK, D_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSI_nSN_SDFCHK, D_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_nSI_nSN_SDFCHK, nD_nSI_nSN, 1'b1);
    tsmc_xbuf (D_SE_SN_SDFCHK, D_SE_SN, 1'b1);
    tsmc_xbuf (D_SE_nSN_SDFCHK, D_SE_nSN, 1'b1);
    tsmc_xbuf (nD_SE_SN_SDFCHK, nD_SE_SN, 1'b1);
    tsmc_xbuf (nD_SE_nSN_SDFCHK, nD_SE_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nSN, SN);
    and (D_SE_SI_SN, D, SE, SI, SN);
    and (D_SE_SI_nSN, D, SE, SI, nSN);
    and (D_nSE_SI_SN, D, nSE, SI, SN);
    and (D_nSE_SI_nSN, D, nSE, SI, nSN);
    and (D_nSE_nSI_SN, D, nSE, nSI, SN);
    and (D_nSE_nSI_nSN, D, nSE, nSI, nSN);
    and (nD_SE_SI_SN, nD, SE, SI, SN);
    and (nD_SE_SI_nSN, nD, SE, SI, nSN);
    and (nD_nSE_SI_nSN, nD, nSE, SI, nSN);
    and (nD_nSE_nSI_nSN, nD, nSE, nSI, nSN);
    and (D_SE_nSI_SN, D, SE, nSI, SN);
    and (D_SE_nSI_nSN, D, SE, nSI, nSN);
    and (nD_SE_nSI_SN, nD, SE, nSI, SN);
    and (nD_SE_nSI_nSN, nD, SE, nSI, nSN);
    and (nD_nSE_SI_SN, nD, nSE, SI, SN);
    and (nD_nSE_nSI_SN, nD, nSE, nSI, SN);
    and (nSE_SI_SN, nSE, SI, SN);
    and (nSE_nSI_SN, nSE, nSI, SN);
    and (nD_SI_SN, nD, SI, SN);
    and (D_nSI_SN, D, nSI, SN);
    and (D_nSI_nSN, D, nSI, nSN);
    and (nD_nSI_nSN, nD, nSI, nSN);
    and (D_SE_SN, D, SE, SN);
    and (D_SE_nSN, D, SE, nSN);
    and (nD_SE_SN, nD, SE, SN);
    and (nD_SE_nSN, nD, SE, nSN);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, SN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, SN);
  `endif
  buf  (SN_check, SE_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKSNQD4 (SI, D, SE, CP, SN, Q);
    input SI, D, SE, CP, SN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (D1, S, D_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (D1, S, D);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SN_SDFCHK, D_SE_SI_SN, 1'b1);
    tsmc_xbuf (D_SE_SI_nSN_SDFCHK, D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_SI_SN_SDFCHK, D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (D_nSE_SI_nSN_SDFCHK, D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SN_SDFCHK, D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_nSN_SDFCHK, D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_SE_SI_SN_SDFCHK, nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (nD_SE_SI_nSN_SDFCHK, nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_nSN_SDFCHK, nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_nSN_SDFCHK, nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (D_SE_nSI_SN_SDFCHK, D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (D_SE_nSI_nSN_SDFCHK, D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SN_SDFCHK, nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nD_SE_nSI_nSN_SDFCHK, nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SN_SDFCHK, nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SN_SDFCHK, nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nSE_SI_SN_SDFCHK, nSE_SI_SN, 1'b1);
    tsmc_xbuf (nSE_nSI_SN_SDFCHK, nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nD_SI_SN_SDFCHK, nD_SI_SN, 1'b1);
    tsmc_xbuf (D_nSI_SN_SDFCHK, D_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSI_nSN_SDFCHK, D_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_nSI_nSN_SDFCHK, nD_nSI_nSN, 1'b1);
    tsmc_xbuf (D_SE_SN_SDFCHK, D_SE_SN, 1'b1);
    tsmc_xbuf (D_SE_nSN_SDFCHK, D_SE_nSN, 1'b1);
    tsmc_xbuf (nD_SE_SN_SDFCHK, nD_SE_SN, 1'b1);
    tsmc_xbuf (nD_SE_nSN_SDFCHK, nD_SE_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nSN, SN);
    and (D_SE_SI_SN, D, SE, SI, SN);
    and (D_SE_SI_nSN, D, SE, SI, nSN);
    and (D_nSE_SI_SN, D, nSE, SI, SN);
    and (D_nSE_SI_nSN, D, nSE, SI, nSN);
    and (D_nSE_nSI_SN, D, nSE, nSI, SN);
    and (D_nSE_nSI_nSN, D, nSE, nSI, nSN);
    and (nD_SE_SI_SN, nD, SE, SI, SN);
    and (nD_SE_SI_nSN, nD, SE, SI, nSN);
    and (nD_nSE_SI_nSN, nD, nSE, SI, nSN);
    and (nD_nSE_nSI_nSN, nD, nSE, nSI, nSN);
    and (D_SE_nSI_SN, D, SE, nSI, SN);
    and (D_SE_nSI_nSN, D, SE, nSI, nSN);
    and (nD_SE_nSI_SN, nD, SE, nSI, SN);
    and (nD_SE_nSI_nSN, nD, SE, nSI, nSN);
    and (nD_nSE_SI_SN, nD, nSE, SI, SN);
    and (nD_nSE_nSI_SN, nD, nSE, nSI, SN);
    and (nSE_SI_SN, nSE, SI, SN);
    and (nSE_nSI_SN, nSE, nSI, SN);
    and (nD_SI_SN, nD, SI, SN);
    and (D_nSI_SN, D, nSI, SN);
    and (D_nSI_nSN, D, nSI, nSN);
    and (nD_nSI_nSN, nD, nSI, nSN);
    and (D_SE_SN, D, SE, SN);
    and (D_SE_nSN, D, SE, nSN);
    and (nD_SE_SN, nD, SE, SN);
    and (nD_SE_nSN, nD, SE, nSN);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, SN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, SN);
  `endif
  buf  (SN_check, SE_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNCND0 (SI, D, SE, CPN, CDN, Q, QN);
    input SI, D, SE, CPN, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CPN_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_D_SE_SI_SDFCHK, CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SE_nSI_SDFCHK, CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_SI_SDFCHK, CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_nSI_SDFCHK, CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_SI_SDFCHK, CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_nSI_SDFCHK, CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_SI_SDFCHK, CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_nSI_SDFCHK, CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_SI_SDFCHK, nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_nSI_SDFCHK, nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_SI_SDFCHK, nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_nSI_SDFCHK, nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_SI_SDFCHK, nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_nSI_SDFCHK, nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_SI_SDFCHK, nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_nSI_SDFCHK, nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCPN, CPN);
    and (CPN_D_SE_SI, CPN, D, SE, SI);
    and (CPN_D_SE_nSI, CPN, D, SE, nSI);
    and (CPN_D_nSE_SI, CPN, D, nSE, SI);
    and (CPN_D_nSE_nSI, CPN, D, nSE, nSI);
    and (CPN_nD_SE_SI, CPN, nD, SE, SI);
    and (CPN_nD_SE_nSI, CPN, nD, SE, nSI);
    and (CPN_nD_nSE_SI, CPN, nD, nSE, SI);
    and (CPN_nD_nSE_nSI, CPN, nD, nSE, nSI);
    and (nCPN_D_SE_SI, nCPN, D, SE, SI);
    and (nCPN_D_SE_nSI, nCPN, D, SE, nSI);
    and (nCPN_D_nSE_SI, nCPN, D, nSE, SI);
    and (nCPN_D_nSE_nSI, nCPN, D, nSE, nSI);
    and (nCPN_nD_SE_SI, nCPN, nD, SE, SI);
    and (nCPN_nD_SE_nSI, nCPN, nD, SE, nSI);
    and (nCPN_nD_nSE_SI, nCPN, nD, nSE, SI);
    and (nCPN_nD_nSE_nSI, nCPN, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
  `endif
  and  (D_check, CDN_i, SE_int_not);
  buf  (CPN_check, CDN_i);
  buf  (SE_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, negedge CPN &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, negedge CPN &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, negedge CPN &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, negedge CPN &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, negedge CPN &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, negedge CPN &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, negedge CPN &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, negedge CPN &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, negedge CPN &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, negedge CPN &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, negedge CPN &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, negedge CPN &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNCND1 (SI, D, SE, CPN, CDN, Q, QN);
    input SI, D, SE, CPN, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CPN_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_D_SE_SI_SDFCHK, CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SE_nSI_SDFCHK, CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_SI_SDFCHK, CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_nSI_SDFCHK, CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_SI_SDFCHK, CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_nSI_SDFCHK, CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_SI_SDFCHK, CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_nSI_SDFCHK, CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_SI_SDFCHK, nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_nSI_SDFCHK, nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_SI_SDFCHK, nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_nSI_SDFCHK, nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_SI_SDFCHK, nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_nSI_SDFCHK, nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_SI_SDFCHK, nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_nSI_SDFCHK, nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCPN, CPN);
    and (CPN_D_SE_SI, CPN, D, SE, SI);
    and (CPN_D_SE_nSI, CPN, D, SE, nSI);
    and (CPN_D_nSE_SI, CPN, D, nSE, SI);
    and (CPN_D_nSE_nSI, CPN, D, nSE, nSI);
    and (CPN_nD_SE_SI, CPN, nD, SE, SI);
    and (CPN_nD_SE_nSI, CPN, nD, SE, nSI);
    and (CPN_nD_nSE_SI, CPN, nD, nSE, SI);
    and (CPN_nD_nSE_nSI, CPN, nD, nSE, nSI);
    and (nCPN_D_SE_SI, nCPN, D, SE, SI);
    and (nCPN_D_SE_nSI, nCPN, D, SE, nSI);
    and (nCPN_D_nSE_SI, nCPN, D, nSE, SI);
    and (nCPN_D_nSE_nSI, nCPN, D, nSE, nSI);
    and (nCPN_nD_SE_SI, nCPN, nD, SE, SI);
    and (nCPN_nD_SE_nSI, nCPN, nD, SE, nSI);
    and (nCPN_nD_nSE_SI, nCPN, nD, nSE, SI);
    and (nCPN_nD_nSE_nSI, nCPN, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
  `endif
  and  (D_check, CDN_i, SE_int_not);
  buf  (CPN_check, CDN_i);
  buf  (SE_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, negedge CPN &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, negedge CPN &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, negedge CPN &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, negedge CPN &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, negedge CPN &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, negedge CPN &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, negedge CPN &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, negedge CPN &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, negedge CPN &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, negedge CPN &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, negedge CPN &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, negedge CPN &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNCND2 (SI, D, SE, CPN, CDN, Q, QN);
    input SI, D, SE, CPN, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CPN_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_D_SE_SI_SDFCHK, CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SE_nSI_SDFCHK, CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_SI_SDFCHK, CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_nSI_SDFCHK, CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_SI_SDFCHK, CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_nSI_SDFCHK, CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_SI_SDFCHK, CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_nSI_SDFCHK, CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_SI_SDFCHK, nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_nSI_SDFCHK, nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_SI_SDFCHK, nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_nSI_SDFCHK, nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_SI_SDFCHK, nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_nSI_SDFCHK, nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_SI_SDFCHK, nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_nSI_SDFCHK, nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCPN, CPN);
    and (CPN_D_SE_SI, CPN, D, SE, SI);
    and (CPN_D_SE_nSI, CPN, D, SE, nSI);
    and (CPN_D_nSE_SI, CPN, D, nSE, SI);
    and (CPN_D_nSE_nSI, CPN, D, nSE, nSI);
    and (CPN_nD_SE_SI, CPN, nD, SE, SI);
    and (CPN_nD_SE_nSI, CPN, nD, SE, nSI);
    and (CPN_nD_nSE_SI, CPN, nD, nSE, SI);
    and (CPN_nD_nSE_nSI, CPN, nD, nSE, nSI);
    and (nCPN_D_SE_SI, nCPN, D, SE, SI);
    and (nCPN_D_SE_nSI, nCPN, D, SE, nSI);
    and (nCPN_D_nSE_SI, nCPN, D, nSE, SI);
    and (nCPN_D_nSE_nSI, nCPN, D, nSE, nSI);
    and (nCPN_nD_SE_SI, nCPN, nD, SE, SI);
    and (nCPN_nD_SE_nSI, nCPN, nD, SE, nSI);
    and (nCPN_nD_nSE_SI, nCPN, nD, nSE, SI);
    and (nCPN_nD_nSE_nSI, nCPN, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
  `endif
  and  (D_check, CDN_i, SE_int_not);
  buf  (CPN_check, CDN_i);
  buf  (SE_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, negedge CPN &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, negedge CPN &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, negedge CPN &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, negedge CPN &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, negedge CPN &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, negedge CPN &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, negedge CPN &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, negedge CPN &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, negedge CPN &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, negedge CPN &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, negedge CPN &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, negedge CPN &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNCND4 (SI, D, SE, CPN, CDN, Q, QN);
    input SI, D, SE, CPN, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CPN_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_D_SE_SI_SDFCHK, CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SE_nSI_SDFCHK, CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_SI_SDFCHK, CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_nSI_SDFCHK, CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_SI_SDFCHK, CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_nSI_SDFCHK, CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_SI_SDFCHK, CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_nSI_SDFCHK, CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_SI_SDFCHK, nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_nSI_SDFCHK, nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_SI_SDFCHK, nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_nSI_SDFCHK, nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_SI_SDFCHK, nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_nSI_SDFCHK, nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_SI_SDFCHK, nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_nSI_SDFCHK, nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCPN, CPN);
    and (CPN_D_SE_SI, CPN, D, SE, SI);
    and (CPN_D_SE_nSI, CPN, D, SE, nSI);
    and (CPN_D_nSE_SI, CPN, D, nSE, SI);
    and (CPN_D_nSE_nSI, CPN, D, nSE, nSI);
    and (CPN_nD_SE_SI, CPN, nD, SE, SI);
    and (CPN_nD_SE_nSI, CPN, nD, SE, nSI);
    and (CPN_nD_nSE_SI, CPN, nD, nSE, SI);
    and (CPN_nD_nSE_nSI, CPN, nD, nSE, nSI);
    and (nCPN_D_SE_SI, nCPN, D, SE, SI);
    and (nCPN_D_SE_nSI, nCPN, D, SE, nSI);
    and (nCPN_D_nSE_SI, nCPN, D, nSE, SI);
    and (nCPN_D_nSE_nSI, nCPN, D, nSE, nSI);
    and (nCPN_nD_SE_SI, nCPN, nD, SE, SI);
    and (nCPN_nD_SE_nSI, nCPN, nD, SE, nSI);
    and (nCPN_nD_nSE_SI, nCPN, nD, nSE, SI);
    and (nCPN_nD_nSE_nSI, nCPN, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
  `endif
  and  (D_check, CDN_i, SE_int_not);
  buf  (CPN_check, CDN_i);
  buf  (SE_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, negedge CPN &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, negedge CPN &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, negedge CPN &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, negedge CPN &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, negedge CPN &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, negedge CPN &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, negedge CPN &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, negedge CPN &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, negedge CPN &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, negedge CPN &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, negedge CPN &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, negedge CPN &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNCSND0 (SI, D, SE, CPN, CDN, SDN, Q, QN);
    input SI, D, SE, CPN, CDN, SDN;
    output Q, QN;
    reg notifier;
    reg flag;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CPN_d;
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_D_SDN_SE_SI_SDFCHK, CPN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SDN_SE_nSI_SDFCHK, CPN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_SDN_nSE_SI_SDFCHK, CPN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SDN_nSE_nSI_SDFCHK, CPN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_SE_SI_SDFCHK, CPN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_SE_nSI_SDFCHK, CPN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_nSE_SI_SDFCHK, CPN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_nSE_nSI_SDFCHK, CPN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_SE_SI_SDFCHK, nCPN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_SE_nSI_SDFCHK, nCPN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_nSE_SI_SDFCHK, nCPN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_nSE_nSI_SDFCHK, nCPN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_SE_SI_SDFCHK, nCPN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_SE_nSI_SDFCHK, nCPN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_nSE_SI_SDFCHK, nCPN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_nSE_nSI_SDFCHK, nCPN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SI_SDFCHK, CDN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_SI_SDFCHK, CDN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_nSI_SDFCHK, CDN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SI_SDFCHK, CDN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_nSI_SDFCHK, CDN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_nSI_SDFCHK, CDN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_SI_SDFCHK, CDN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_nSI_SDFCHK, CDN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_SE_SI_SDFCHK, CDN_CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_nSE_SI_SDFCHK, CDN_CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_nSE_nSI_SDFCHK, CDN_CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_SE_SI_SDFCHK, CDN_CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_SE_nSI_SDFCHK, CDN_CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_SE_nSI_SDFCHK, CDN_CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_nSE_SI_SDFCHK, CDN_CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_nSE_nSI_SDFCHK, CDN_CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_SE_SI_SDFCHK, CDN_nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_SE_nSI_SDFCHK, CDN_nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_nSE_SI_SDFCHK, CDN_nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_nSE_nSI_SDFCHK, CDN_nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_SE_SI_SDFCHK, CDN_nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_SE_nSI_SDFCHK, CDN_nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_nSE_SI_SDFCHK, CDN_nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_nSE_nSI_SDFCHK, CDN_nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_SE_SI_SDFCHK, CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_SI_SDFCHK, CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_nSI_SDFCHK, CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_SI_SDFCHK, CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SE_nSI_SDFCHK, CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_nSI_SDFCHK, CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_SI_SDFCHK, CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_nSI_SDFCHK, CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_SI_SDFCHK, nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_nSI_SDFCHK, nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_SI_SDFCHK, nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_nSI_SDFCHK, nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_SI_SDFCHK, nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_nSI_SDFCHK, nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_SI_SDFCHK, nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_nSI_SDFCHK, nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_SI_SDFCHK, CDN_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_nSI_SDFCHK, CDN_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SI_SDFCHK, CDN_nD_SDN_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSI_SDFCHK, CDN_D_SDN_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SDFCHK, CDN_D_SDN_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SDFCHK, CDN_nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCPN, CPN);
    and (CPN_D_SDN_SE_SI, CPN, D, SDN, SE, SI);
    and (CPN_D_SDN_SE_nSI, CPN, D, SDN, SE, nSI);
    and (CPN_D_SDN_nSE_SI, CPN, D, SDN, nSE, SI);
    and (CPN_D_SDN_nSE_nSI, CPN, D, SDN, nSE, nSI);
    and (CPN_nD_SDN_SE_SI, CPN, nD, SDN, SE, SI);
    and (CPN_nD_SDN_SE_nSI, CPN, nD, SDN, SE, nSI);
    and (CPN_nD_SDN_nSE_SI, CPN, nD, SDN, nSE, SI);
    and (CPN_nD_SDN_nSE_nSI, CPN, nD, SDN, nSE, nSI);
    and (nCPN_D_SDN_SE_SI, nCPN, D, SDN, SE, SI);
    and (nCPN_D_SDN_SE_nSI, nCPN, D, SDN, SE, nSI);
    and (nCPN_D_SDN_nSE_SI, nCPN, D, SDN, nSE, SI);
    and (nCPN_D_SDN_nSE_nSI, nCPN, D, SDN, nSE, nSI);
    and (nCPN_nD_SDN_SE_SI, nCPN, nD, SDN, SE, SI);
    and (nCPN_nD_SDN_SE_nSI, nCPN, nD, SDN, SE, nSI);
    and (nCPN_nD_SDN_nSE_SI, nCPN, nD, SDN, nSE, SI);
    and (nCPN_nD_SDN_nSE_nSI, nCPN, nD, SDN, nSE, nSI);
    and (CDN_D_SDN_SE_SI, CDN, D, SDN, SE, SI);
    and (CDN_D_SDN_nSE_SI, CDN, D, SDN, nSE, SI);
    and (CDN_D_SDN_nSE_nSI, CDN, D, SDN, nSE, nSI);
    and (CDN_nD_SDN_SE_SI, CDN, nD, SDN, SE, SI);
    and (CDN_D_SDN_SE_nSI, CDN, D, SDN, SE, nSI);
    and (CDN_nD_SDN_SE_nSI, CDN, nD, SDN, SE, nSI);
    and (CDN_nD_SDN_nSE_SI, CDN, nD, SDN, nSE, SI);
    and (CDN_nD_SDN_nSE_nSI, CDN, nD, SDN, nSE, nSI);
    and (CDN_CPN_D_SE_SI, CDN, CPN, D, SE, SI);
    and (CDN_CPN_D_nSE_SI, CDN, CPN, D, nSE, SI);
    and (CDN_CPN_D_nSE_nSI, CDN, CPN, D, nSE, nSI);
    and (CDN_CPN_nD_SE_SI, CDN, CPN, nD, SE, SI);
    and (CDN_CPN_D_SE_nSI, CDN, CPN, D, SE, nSI);
    and (CDN_CPN_nD_SE_nSI, CDN, CPN, nD, SE, nSI);
    and (CDN_CPN_nD_nSE_SI, CDN, CPN, nD, nSE, SI);
    and (CDN_CPN_nD_nSE_nSI, CDN, CPN, nD, nSE, nSI);
    and (CDN_nCPN_D_SE_SI, CDN, nCPN, D, SE, SI);
    and (CDN_nCPN_D_SE_nSI, CDN, nCPN, D, SE, nSI);
    and (CDN_nCPN_D_nSE_SI, CDN, nCPN, D, nSE, SI);
    and (CDN_nCPN_D_nSE_nSI, CDN, nCPN, D, nSE, nSI);
    and (CDN_nCPN_nD_SE_SI, CDN, nCPN, nD, SE, SI);
    and (CDN_nCPN_nD_SE_nSI, CDN, nCPN, nD, SE, nSI);
    and (CDN_nCPN_nD_nSE_SI, CDN, nCPN, nD, nSE, SI);
    and (CDN_nCPN_nD_nSE_nSI, CDN, nCPN, nD, nSE, nSI);
    and (CPN_D_SE_SI, CPN, D, SE, SI);
    and (CPN_D_nSE_SI, CPN, D, nSE, SI);
    and (CPN_D_nSE_nSI, CPN, D, nSE, nSI);
    and (CPN_nD_SE_SI, CPN, nD, SE, SI);
    and (CPN_D_SE_nSI, CPN, D, SE, nSI);
    and (CPN_nD_SE_nSI, CPN, nD, SE, nSI);
    and (CPN_nD_nSE_SI, CPN, nD, nSE, SI);
    and (CPN_nD_nSE_nSI, CPN, nD, nSE, nSI);
    and (nCPN_D_SE_SI, nCPN, D, SE, SI);
    and (nCPN_D_SE_nSI, nCPN, D, SE, nSI);
    and (nCPN_D_nSE_SI, nCPN, D, nSE, SI);
    and (nCPN_D_nSE_nSI, nCPN, D, nSE, nSI);
    and (nCPN_nD_SE_SI, nCPN, nD, SE, SI);
    and (nCPN_nD_SE_nSI, nCPN, nD, SE, nSI);
    and (nCPN_nD_nSE_SI, nCPN, nD, nSE, SI);
    and (nCPN_nD_nSE_nSI, nCPN, nD, nSE, nSI);
    and (CDN_SDN_nSE_SI, CDN, SDN, nSE, SI);
    and (CDN_SDN_nSE_nSI, CDN, SDN, nSE, nSI);
    and (CDN_nD_SDN_SI, CDN, nD, SDN, SI);
    and (CDN_D_SDN_nSI, CDN, D, SDN, nSI);
    and (CDN_D_SDN_SE, CDN, D, SDN, SE);
    and (CDN_nD_SDN_SE, CDN, nD, SDN, SE);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SDN_i, SE);
  `endif
  and  (D_check, CDN_i, SDN_i, SE_int_not);
  and  (CPN_check, CDN_i, SDN_i);
  and  (SE_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge CDN &&& CPN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (posedge CDN &&& CPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge CDN &&& D_SDN_SE_SI_SDFCHK, negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (posedge SDN &&& CPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (posedge CDN &&& CPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNCSND1 (SI, D, SE, CPN, CDN, SDN, Q, QN);
    input SI, D, SE, CPN, CDN, SDN;
    output Q, QN;
    reg notifier;
    reg flag;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CPN_d;
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_D_SDN_SE_SI_SDFCHK, CPN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SDN_SE_nSI_SDFCHK, CPN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_SDN_nSE_SI_SDFCHK, CPN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SDN_nSE_nSI_SDFCHK, CPN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_SE_SI_SDFCHK, CPN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_SE_nSI_SDFCHK, CPN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_nSE_SI_SDFCHK, CPN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_nSE_nSI_SDFCHK, CPN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_SE_SI_SDFCHK, nCPN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_SE_nSI_SDFCHK, nCPN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_nSE_SI_SDFCHK, nCPN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_nSE_nSI_SDFCHK, nCPN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_SE_SI_SDFCHK, nCPN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_SE_nSI_SDFCHK, nCPN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_nSE_SI_SDFCHK, nCPN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_nSE_nSI_SDFCHK, nCPN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SI_SDFCHK, CDN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_SI_SDFCHK, CDN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_nSI_SDFCHK, CDN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SI_SDFCHK, CDN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_nSI_SDFCHK, CDN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_nSI_SDFCHK, CDN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_SI_SDFCHK, CDN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_nSI_SDFCHK, CDN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_SE_SI_SDFCHK, CDN_CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_nSE_SI_SDFCHK, CDN_CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_nSE_nSI_SDFCHK, CDN_CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_SE_SI_SDFCHK, CDN_CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_SE_nSI_SDFCHK, CDN_CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_SE_nSI_SDFCHK, CDN_CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_nSE_SI_SDFCHK, CDN_CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_nSE_nSI_SDFCHK, CDN_CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_SE_SI_SDFCHK, CDN_nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_SE_nSI_SDFCHK, CDN_nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_nSE_SI_SDFCHK, CDN_nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_nSE_nSI_SDFCHK, CDN_nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_SE_SI_SDFCHK, CDN_nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_SE_nSI_SDFCHK, CDN_nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_nSE_SI_SDFCHK, CDN_nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_nSE_nSI_SDFCHK, CDN_nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_SE_SI_SDFCHK, CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_SI_SDFCHK, CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_nSI_SDFCHK, CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_SI_SDFCHK, CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SE_nSI_SDFCHK, CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_nSI_SDFCHK, CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_SI_SDFCHK, CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_nSI_SDFCHK, CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_SI_SDFCHK, nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_nSI_SDFCHK, nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_SI_SDFCHK, nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_nSI_SDFCHK, nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_SI_SDFCHK, nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_nSI_SDFCHK, nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_SI_SDFCHK, nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_nSI_SDFCHK, nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_SI_SDFCHK, CDN_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_nSI_SDFCHK, CDN_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SI_SDFCHK, CDN_nD_SDN_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSI_SDFCHK, CDN_D_SDN_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SDFCHK, CDN_D_SDN_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SDFCHK, CDN_nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCPN, CPN);
    and (CPN_D_SDN_SE_SI, CPN, D, SDN, SE, SI);
    and (CPN_D_SDN_SE_nSI, CPN, D, SDN, SE, nSI);
    and (CPN_D_SDN_nSE_SI, CPN, D, SDN, nSE, SI);
    and (CPN_D_SDN_nSE_nSI, CPN, D, SDN, nSE, nSI);
    and (CPN_nD_SDN_SE_SI, CPN, nD, SDN, SE, SI);
    and (CPN_nD_SDN_SE_nSI, CPN, nD, SDN, SE, nSI);
    and (CPN_nD_SDN_nSE_SI, CPN, nD, SDN, nSE, SI);
    and (CPN_nD_SDN_nSE_nSI, CPN, nD, SDN, nSE, nSI);
    and (nCPN_D_SDN_SE_SI, nCPN, D, SDN, SE, SI);
    and (nCPN_D_SDN_SE_nSI, nCPN, D, SDN, SE, nSI);
    and (nCPN_D_SDN_nSE_SI, nCPN, D, SDN, nSE, SI);
    and (nCPN_D_SDN_nSE_nSI, nCPN, D, SDN, nSE, nSI);
    and (nCPN_nD_SDN_SE_SI, nCPN, nD, SDN, SE, SI);
    and (nCPN_nD_SDN_SE_nSI, nCPN, nD, SDN, SE, nSI);
    and (nCPN_nD_SDN_nSE_SI, nCPN, nD, SDN, nSE, SI);
    and (nCPN_nD_SDN_nSE_nSI, nCPN, nD, SDN, nSE, nSI);
    and (CDN_D_SDN_SE_SI, CDN, D, SDN, SE, SI);
    and (CDN_D_SDN_nSE_SI, CDN, D, SDN, nSE, SI);
    and (CDN_D_SDN_nSE_nSI, CDN, D, SDN, nSE, nSI);
    and (CDN_nD_SDN_SE_SI, CDN, nD, SDN, SE, SI);
    and (CDN_D_SDN_SE_nSI, CDN, D, SDN, SE, nSI);
    and (CDN_nD_SDN_SE_nSI, CDN, nD, SDN, SE, nSI);
    and (CDN_nD_SDN_nSE_SI, CDN, nD, SDN, nSE, SI);
    and (CDN_nD_SDN_nSE_nSI, CDN, nD, SDN, nSE, nSI);
    and (CDN_CPN_D_SE_SI, CDN, CPN, D, SE, SI);
    and (CDN_CPN_D_nSE_SI, CDN, CPN, D, nSE, SI);
    and (CDN_CPN_D_nSE_nSI, CDN, CPN, D, nSE, nSI);
    and (CDN_CPN_nD_SE_SI, CDN, CPN, nD, SE, SI);
    and (CDN_CPN_D_SE_nSI, CDN, CPN, D, SE, nSI);
    and (CDN_CPN_nD_SE_nSI, CDN, CPN, nD, SE, nSI);
    and (CDN_CPN_nD_nSE_SI, CDN, CPN, nD, nSE, SI);
    and (CDN_CPN_nD_nSE_nSI, CDN, CPN, nD, nSE, nSI);
    and (CDN_nCPN_D_SE_SI, CDN, nCPN, D, SE, SI);
    and (CDN_nCPN_D_SE_nSI, CDN, nCPN, D, SE, nSI);
    and (CDN_nCPN_D_nSE_SI, CDN, nCPN, D, nSE, SI);
    and (CDN_nCPN_D_nSE_nSI, CDN, nCPN, D, nSE, nSI);
    and (CDN_nCPN_nD_SE_SI, CDN, nCPN, nD, SE, SI);
    and (CDN_nCPN_nD_SE_nSI, CDN, nCPN, nD, SE, nSI);
    and (CDN_nCPN_nD_nSE_SI, CDN, nCPN, nD, nSE, SI);
    and (CDN_nCPN_nD_nSE_nSI, CDN, nCPN, nD, nSE, nSI);
    and (CPN_D_SE_SI, CPN, D, SE, SI);
    and (CPN_D_nSE_SI, CPN, D, nSE, SI);
    and (CPN_D_nSE_nSI, CPN, D, nSE, nSI);
    and (CPN_nD_SE_SI, CPN, nD, SE, SI);
    and (CPN_D_SE_nSI, CPN, D, SE, nSI);
    and (CPN_nD_SE_nSI, CPN, nD, SE, nSI);
    and (CPN_nD_nSE_SI, CPN, nD, nSE, SI);
    and (CPN_nD_nSE_nSI, CPN, nD, nSE, nSI);
    and (nCPN_D_SE_SI, nCPN, D, SE, SI);
    and (nCPN_D_SE_nSI, nCPN, D, SE, nSI);
    and (nCPN_D_nSE_SI, nCPN, D, nSE, SI);
    and (nCPN_D_nSE_nSI, nCPN, D, nSE, nSI);
    and (nCPN_nD_SE_SI, nCPN, nD, SE, SI);
    and (nCPN_nD_SE_nSI, nCPN, nD, SE, nSI);
    and (nCPN_nD_nSE_SI, nCPN, nD, nSE, SI);
    and (nCPN_nD_nSE_nSI, nCPN, nD, nSE, nSI);
    and (CDN_SDN_nSE_SI, CDN, SDN, nSE, SI);
    and (CDN_SDN_nSE_nSI, CDN, SDN, nSE, nSI);
    and (CDN_nD_SDN_SI, CDN, nD, SDN, SI);
    and (CDN_D_SDN_nSI, CDN, D, SDN, nSI);
    and (CDN_D_SDN_SE, CDN, D, SDN, SE);
    and (CDN_nD_SDN_SE, CDN, nD, SDN, SE);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SDN_i, SE);
  `endif
  and  (D_check, CDN_i, SDN_i, SE_int_not);
  and  (CPN_check, CDN_i, SDN_i);
  and  (SE_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge CDN &&& CPN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (posedge CDN &&& CPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge CDN &&& D_SDN_SE_SI_SDFCHK, negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (posedge SDN &&& CPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (posedge CDN &&& CPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNCSND2 (SI, D, SE, CPN, CDN, SDN, Q, QN);
    input SI, D, SE, CPN, CDN, SDN;
    output Q, QN;
    reg notifier;
    reg flag;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CPN_d;
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_D_SDN_SE_SI_SDFCHK, CPN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SDN_SE_nSI_SDFCHK, CPN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_SDN_nSE_SI_SDFCHK, CPN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SDN_nSE_nSI_SDFCHK, CPN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_SE_SI_SDFCHK, CPN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_SE_nSI_SDFCHK, CPN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_nSE_SI_SDFCHK, CPN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_nSE_nSI_SDFCHK, CPN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_SE_SI_SDFCHK, nCPN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_SE_nSI_SDFCHK, nCPN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_nSE_SI_SDFCHK, nCPN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_nSE_nSI_SDFCHK, nCPN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_SE_SI_SDFCHK, nCPN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_SE_nSI_SDFCHK, nCPN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_nSE_SI_SDFCHK, nCPN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_nSE_nSI_SDFCHK, nCPN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SI_SDFCHK, CDN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_SI_SDFCHK, CDN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_nSI_SDFCHK, CDN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SI_SDFCHK, CDN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_nSI_SDFCHK, CDN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_nSI_SDFCHK, CDN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_SI_SDFCHK, CDN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_nSI_SDFCHK, CDN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_SE_SI_SDFCHK, CDN_CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_nSE_SI_SDFCHK, CDN_CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_nSE_nSI_SDFCHK, CDN_CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_SE_SI_SDFCHK, CDN_CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_SE_nSI_SDFCHK, CDN_CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_SE_nSI_SDFCHK, CDN_CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_nSE_SI_SDFCHK, CDN_CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_nSE_nSI_SDFCHK, CDN_CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_SE_SI_SDFCHK, CDN_nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_SE_nSI_SDFCHK, CDN_nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_nSE_SI_SDFCHK, CDN_nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_nSE_nSI_SDFCHK, CDN_nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_SE_SI_SDFCHK, CDN_nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_SE_nSI_SDFCHK, CDN_nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_nSE_SI_SDFCHK, CDN_nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_nSE_nSI_SDFCHK, CDN_nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_SE_SI_SDFCHK, CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_SI_SDFCHK, CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_nSI_SDFCHK, CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_SI_SDFCHK, CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SE_nSI_SDFCHK, CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_nSI_SDFCHK, CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_SI_SDFCHK, CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_nSI_SDFCHK, CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_SI_SDFCHK, nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_nSI_SDFCHK, nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_SI_SDFCHK, nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_nSI_SDFCHK, nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_SI_SDFCHK, nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_nSI_SDFCHK, nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_SI_SDFCHK, nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_nSI_SDFCHK, nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_SI_SDFCHK, CDN_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_nSI_SDFCHK, CDN_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SI_SDFCHK, CDN_nD_SDN_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSI_SDFCHK, CDN_D_SDN_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SDFCHK, CDN_D_SDN_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SDFCHK, CDN_nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCPN, CPN);
    and (CPN_D_SDN_SE_SI, CPN, D, SDN, SE, SI);
    and (CPN_D_SDN_SE_nSI, CPN, D, SDN, SE, nSI);
    and (CPN_D_SDN_nSE_SI, CPN, D, SDN, nSE, SI);
    and (CPN_D_SDN_nSE_nSI, CPN, D, SDN, nSE, nSI);
    and (CPN_nD_SDN_SE_SI, CPN, nD, SDN, SE, SI);
    and (CPN_nD_SDN_SE_nSI, CPN, nD, SDN, SE, nSI);
    and (CPN_nD_SDN_nSE_SI, CPN, nD, SDN, nSE, SI);
    and (CPN_nD_SDN_nSE_nSI, CPN, nD, SDN, nSE, nSI);
    and (nCPN_D_SDN_SE_SI, nCPN, D, SDN, SE, SI);
    and (nCPN_D_SDN_SE_nSI, nCPN, D, SDN, SE, nSI);
    and (nCPN_D_SDN_nSE_SI, nCPN, D, SDN, nSE, SI);
    and (nCPN_D_SDN_nSE_nSI, nCPN, D, SDN, nSE, nSI);
    and (nCPN_nD_SDN_SE_SI, nCPN, nD, SDN, SE, SI);
    and (nCPN_nD_SDN_SE_nSI, nCPN, nD, SDN, SE, nSI);
    and (nCPN_nD_SDN_nSE_SI, nCPN, nD, SDN, nSE, SI);
    and (nCPN_nD_SDN_nSE_nSI, nCPN, nD, SDN, nSE, nSI);
    and (CDN_D_SDN_SE_SI, CDN, D, SDN, SE, SI);
    and (CDN_D_SDN_nSE_SI, CDN, D, SDN, nSE, SI);
    and (CDN_D_SDN_nSE_nSI, CDN, D, SDN, nSE, nSI);
    and (CDN_nD_SDN_SE_SI, CDN, nD, SDN, SE, SI);
    and (CDN_D_SDN_SE_nSI, CDN, D, SDN, SE, nSI);
    and (CDN_nD_SDN_SE_nSI, CDN, nD, SDN, SE, nSI);
    and (CDN_nD_SDN_nSE_SI, CDN, nD, SDN, nSE, SI);
    and (CDN_nD_SDN_nSE_nSI, CDN, nD, SDN, nSE, nSI);
    and (CDN_CPN_D_SE_SI, CDN, CPN, D, SE, SI);
    and (CDN_CPN_D_nSE_SI, CDN, CPN, D, nSE, SI);
    and (CDN_CPN_D_nSE_nSI, CDN, CPN, D, nSE, nSI);
    and (CDN_CPN_nD_SE_SI, CDN, CPN, nD, SE, SI);
    and (CDN_CPN_D_SE_nSI, CDN, CPN, D, SE, nSI);
    and (CDN_CPN_nD_SE_nSI, CDN, CPN, nD, SE, nSI);
    and (CDN_CPN_nD_nSE_SI, CDN, CPN, nD, nSE, SI);
    and (CDN_CPN_nD_nSE_nSI, CDN, CPN, nD, nSE, nSI);
    and (CDN_nCPN_D_SE_SI, CDN, nCPN, D, SE, SI);
    and (CDN_nCPN_D_SE_nSI, CDN, nCPN, D, SE, nSI);
    and (CDN_nCPN_D_nSE_SI, CDN, nCPN, D, nSE, SI);
    and (CDN_nCPN_D_nSE_nSI, CDN, nCPN, D, nSE, nSI);
    and (CDN_nCPN_nD_SE_SI, CDN, nCPN, nD, SE, SI);
    and (CDN_nCPN_nD_SE_nSI, CDN, nCPN, nD, SE, nSI);
    and (CDN_nCPN_nD_nSE_SI, CDN, nCPN, nD, nSE, SI);
    and (CDN_nCPN_nD_nSE_nSI, CDN, nCPN, nD, nSE, nSI);
    and (CPN_D_SE_SI, CPN, D, SE, SI);
    and (CPN_D_nSE_SI, CPN, D, nSE, SI);
    and (CPN_D_nSE_nSI, CPN, D, nSE, nSI);
    and (CPN_nD_SE_SI, CPN, nD, SE, SI);
    and (CPN_D_SE_nSI, CPN, D, SE, nSI);
    and (CPN_nD_SE_nSI, CPN, nD, SE, nSI);
    and (CPN_nD_nSE_SI, CPN, nD, nSE, SI);
    and (CPN_nD_nSE_nSI, CPN, nD, nSE, nSI);
    and (nCPN_D_SE_SI, nCPN, D, SE, SI);
    and (nCPN_D_SE_nSI, nCPN, D, SE, nSI);
    and (nCPN_D_nSE_SI, nCPN, D, nSE, SI);
    and (nCPN_D_nSE_nSI, nCPN, D, nSE, nSI);
    and (nCPN_nD_SE_SI, nCPN, nD, SE, SI);
    and (nCPN_nD_SE_nSI, nCPN, nD, SE, nSI);
    and (nCPN_nD_nSE_SI, nCPN, nD, nSE, SI);
    and (nCPN_nD_nSE_nSI, nCPN, nD, nSE, nSI);
    and (CDN_SDN_nSE_SI, CDN, SDN, nSE, SI);
    and (CDN_SDN_nSE_nSI, CDN, SDN, nSE, nSI);
    and (CDN_nD_SDN_SI, CDN, nD, SDN, SI);
    and (CDN_D_SDN_nSI, CDN, D, SDN, nSI);
    and (CDN_D_SDN_SE, CDN, D, SDN, SE);
    and (CDN_nD_SDN_SE, CDN, nD, SDN, SE);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SDN_i, SE);
  `endif
  and  (D_check, CDN_i, SDN_i, SE_int_not);
  and  (CPN_check, CDN_i, SDN_i);
  and  (SE_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge CDN &&& CPN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (posedge CDN &&& CPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge CDN &&& D_SDN_SE_SI_SDFCHK, negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (posedge SDN &&& CPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (posedge CDN &&& CPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNCSND4 (SI, D, SE, CPN, CDN, SDN, Q, QN);
    input SI, D, SE, CPN, CDN, SDN;
    output Q, QN;
    reg notifier;
    reg flag;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CPN_d;
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_D_SDN_SE_SI_SDFCHK, CPN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SDN_SE_nSI_SDFCHK, CPN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_SDN_nSE_SI_SDFCHK, CPN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SDN_nSE_nSI_SDFCHK, CPN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_SE_SI_SDFCHK, CPN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_SE_nSI_SDFCHK, CPN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_nSE_SI_SDFCHK, CPN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_nSE_nSI_SDFCHK, CPN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_SE_SI_SDFCHK, nCPN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_SE_nSI_SDFCHK, nCPN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_nSE_SI_SDFCHK, nCPN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_nSE_nSI_SDFCHK, nCPN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_SE_SI_SDFCHK, nCPN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_SE_nSI_SDFCHK, nCPN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_nSE_SI_SDFCHK, nCPN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_nSE_nSI_SDFCHK, nCPN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SI_SDFCHK, CDN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_SI_SDFCHK, CDN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_nSI_SDFCHK, CDN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SI_SDFCHK, CDN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_nSI_SDFCHK, CDN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_nSI_SDFCHK, CDN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_SI_SDFCHK, CDN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_nSI_SDFCHK, CDN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_SE_SI_SDFCHK, CDN_CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_nSE_SI_SDFCHK, CDN_CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_nSE_nSI_SDFCHK, CDN_CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_SE_SI_SDFCHK, CDN_CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_SE_nSI_SDFCHK, CDN_CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_SE_nSI_SDFCHK, CDN_CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_nSE_SI_SDFCHK, CDN_CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_nSE_nSI_SDFCHK, CDN_CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_SE_SI_SDFCHK, CDN_nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_SE_nSI_SDFCHK, CDN_nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_nSE_SI_SDFCHK, CDN_nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_nSE_nSI_SDFCHK, CDN_nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_SE_SI_SDFCHK, CDN_nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_SE_nSI_SDFCHK, CDN_nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_nSE_SI_SDFCHK, CDN_nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_nSE_nSI_SDFCHK, CDN_nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_SE_SI_SDFCHK, CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_SI_SDFCHK, CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_nSI_SDFCHK, CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_SI_SDFCHK, CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SE_nSI_SDFCHK, CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_nSI_SDFCHK, CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_SI_SDFCHK, CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_nSI_SDFCHK, CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_SI_SDFCHK, nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_nSI_SDFCHK, nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_SI_SDFCHK, nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_nSI_SDFCHK, nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_SI_SDFCHK, nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_nSI_SDFCHK, nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_SI_SDFCHK, nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_nSI_SDFCHK, nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_SI_SDFCHK, CDN_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_nSI_SDFCHK, CDN_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SI_SDFCHK, CDN_nD_SDN_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSI_SDFCHK, CDN_D_SDN_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SDFCHK, CDN_D_SDN_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SDFCHK, CDN_nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCPN, CPN);
    and (CPN_D_SDN_SE_SI, CPN, D, SDN, SE, SI);
    and (CPN_D_SDN_SE_nSI, CPN, D, SDN, SE, nSI);
    and (CPN_D_SDN_nSE_SI, CPN, D, SDN, nSE, SI);
    and (CPN_D_SDN_nSE_nSI, CPN, D, SDN, nSE, nSI);
    and (CPN_nD_SDN_SE_SI, CPN, nD, SDN, SE, SI);
    and (CPN_nD_SDN_SE_nSI, CPN, nD, SDN, SE, nSI);
    and (CPN_nD_SDN_nSE_SI, CPN, nD, SDN, nSE, SI);
    and (CPN_nD_SDN_nSE_nSI, CPN, nD, SDN, nSE, nSI);
    and (nCPN_D_SDN_SE_SI, nCPN, D, SDN, SE, SI);
    and (nCPN_D_SDN_SE_nSI, nCPN, D, SDN, SE, nSI);
    and (nCPN_D_SDN_nSE_SI, nCPN, D, SDN, nSE, SI);
    and (nCPN_D_SDN_nSE_nSI, nCPN, D, SDN, nSE, nSI);
    and (nCPN_nD_SDN_SE_SI, nCPN, nD, SDN, SE, SI);
    and (nCPN_nD_SDN_SE_nSI, nCPN, nD, SDN, SE, nSI);
    and (nCPN_nD_SDN_nSE_SI, nCPN, nD, SDN, nSE, SI);
    and (nCPN_nD_SDN_nSE_nSI, nCPN, nD, SDN, nSE, nSI);
    and (CDN_D_SDN_SE_SI, CDN, D, SDN, SE, SI);
    and (CDN_D_SDN_nSE_SI, CDN, D, SDN, nSE, SI);
    and (CDN_D_SDN_nSE_nSI, CDN, D, SDN, nSE, nSI);
    and (CDN_nD_SDN_SE_SI, CDN, nD, SDN, SE, SI);
    and (CDN_D_SDN_SE_nSI, CDN, D, SDN, SE, nSI);
    and (CDN_nD_SDN_SE_nSI, CDN, nD, SDN, SE, nSI);
    and (CDN_nD_SDN_nSE_SI, CDN, nD, SDN, nSE, SI);
    and (CDN_nD_SDN_nSE_nSI, CDN, nD, SDN, nSE, nSI);
    and (CDN_CPN_D_SE_SI, CDN, CPN, D, SE, SI);
    and (CDN_CPN_D_nSE_SI, CDN, CPN, D, nSE, SI);
    and (CDN_CPN_D_nSE_nSI, CDN, CPN, D, nSE, nSI);
    and (CDN_CPN_nD_SE_SI, CDN, CPN, nD, SE, SI);
    and (CDN_CPN_D_SE_nSI, CDN, CPN, D, SE, nSI);
    and (CDN_CPN_nD_SE_nSI, CDN, CPN, nD, SE, nSI);
    and (CDN_CPN_nD_nSE_SI, CDN, CPN, nD, nSE, SI);
    and (CDN_CPN_nD_nSE_nSI, CDN, CPN, nD, nSE, nSI);
    and (CDN_nCPN_D_SE_SI, CDN, nCPN, D, SE, SI);
    and (CDN_nCPN_D_SE_nSI, CDN, nCPN, D, SE, nSI);
    and (CDN_nCPN_D_nSE_SI, CDN, nCPN, D, nSE, SI);
    and (CDN_nCPN_D_nSE_nSI, CDN, nCPN, D, nSE, nSI);
    and (CDN_nCPN_nD_SE_SI, CDN, nCPN, nD, SE, SI);
    and (CDN_nCPN_nD_SE_nSI, CDN, nCPN, nD, SE, nSI);
    and (CDN_nCPN_nD_nSE_SI, CDN, nCPN, nD, nSE, SI);
    and (CDN_nCPN_nD_nSE_nSI, CDN, nCPN, nD, nSE, nSI);
    and (CPN_D_SE_SI, CPN, D, SE, SI);
    and (CPN_D_nSE_SI, CPN, D, nSE, SI);
    and (CPN_D_nSE_nSI, CPN, D, nSE, nSI);
    and (CPN_nD_SE_SI, CPN, nD, SE, SI);
    and (CPN_D_SE_nSI, CPN, D, SE, nSI);
    and (CPN_nD_SE_nSI, CPN, nD, SE, nSI);
    and (CPN_nD_nSE_SI, CPN, nD, nSE, SI);
    and (CPN_nD_nSE_nSI, CPN, nD, nSE, nSI);
    and (nCPN_D_SE_SI, nCPN, D, SE, SI);
    and (nCPN_D_SE_nSI, nCPN, D, SE, nSI);
    and (nCPN_D_nSE_SI, nCPN, D, nSE, SI);
    and (nCPN_D_nSE_nSI, nCPN, D, nSE, nSI);
    and (nCPN_nD_SE_SI, nCPN, nD, SE, SI);
    and (nCPN_nD_SE_nSI, nCPN, nD, SE, nSI);
    and (nCPN_nD_nSE_SI, nCPN, nD, nSE, SI);
    and (nCPN_nD_nSE_nSI, nCPN, nD, nSE, nSI);
    and (CDN_SDN_nSE_SI, CDN, SDN, nSE, SI);
    and (CDN_SDN_nSE_nSI, CDN, SDN, nSE, nSI);
    and (CDN_nD_SDN_SI, CDN, nD, SDN, SI);
    and (CDN_D_SDN_nSI, CDN, D, SDN, nSI);
    and (CDN_D_SDN_SE, CDN, D, SDN, SE);
    and (CDN_nD_SDN_SE, CDN, nD, SDN, SE);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SDN_i, SE);
  `endif
  and  (D_check, CDN_i, SDN_i, SE_int_not);
  and  (CPN_check, CDN_i, SDN_i);
  and  (SE_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge CDN &&& CPN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (posedge CDN &&& CPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge CDN &&& D_SDN_SE_SI_SDFCHK, negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (posedge SDN &&& CPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (posedge CDN &&& CPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFND0 (SI, D, SE, CPN, Q, QN);
    input SI, D, SE, CPN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CPN_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CPN_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CPN &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
  `else
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFND1 (SI, D, SE, CPN, Q, QN);
    input SI, D, SE, CPN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CPN_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CPN_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CPN &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
  `else
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFND2 (SI, D, SE, CPN, Q, QN);
    input SI, D, SE, CPN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CPN_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CPN_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CPN &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
  `else
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFND4 (SI, D, SE, CPN, Q, QN);
    input SI, D, SE, CPN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CPN_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CPN_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CPN &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
  `else
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNSND0 (SI, D, SE, CPN, SDN, Q, QN);
    input SI, D, SE, CPN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CPN_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_SE_SI_SDFCHK, CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_SI_SDFCHK, CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_nSI_SDFCHK, CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_SI_SDFCHK, CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SE_nSI_SDFCHK, CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_nSI_SDFCHK, CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_SI_SDFCHK, CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_nSI_SDFCHK, CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_SI_SDFCHK, nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_nSI_SDFCHK, nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_SI_SDFCHK, nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_nSI_SDFCHK, nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_SI_SDFCHK, nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_nSI_SDFCHK, nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_SI_SDFCHK, nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_nSI_SDFCHK, nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCPN, CPN);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CPN_D_SE_SI, CPN, D, SE, SI);
    and (CPN_D_nSE_SI, CPN, D, nSE, SI);
    and (CPN_D_nSE_nSI, CPN, D, nSE, nSI);
    and (CPN_nD_SE_SI, CPN, nD, SE, SI);
    and (CPN_D_SE_nSI, CPN, D, SE, nSI);
    and (CPN_nD_SE_nSI, CPN, nD, SE, nSI);
    and (CPN_nD_nSE_SI, CPN, nD, nSE, SI);
    and (CPN_nD_nSE_nSI, CPN, nD, nSE, nSI);
    and (nCPN_D_SE_SI, nCPN, D, SE, SI);
    and (nCPN_D_SE_nSI, nCPN, D, SE, nSI);
    and (nCPN_D_nSE_SI, nCPN, D, nSE, SI);
    and (nCPN_D_nSE_nSI, nCPN, D, nSE, nSI);
    and (nCPN_nD_SE_SI, nCPN, nD, SE, SI);
    and (nCPN_nD_SE_nSI, nCPN, nD, SE, nSI);
    and (nCPN_nD_nSE_SI, nCPN, nD, nSE, SI);
    and (nCPN_nD_nSE_nSI, nCPN, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, SDN_i, SE);
  `endif
  and  (D_check, SDN_i, SE_int_not);
  buf  (CPN_check, SDN_i);
  buf  (SE_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, negedge CPN &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, negedge CPN &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, negedge CPN &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, negedge CPN &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, negedge CPN &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, negedge CPN &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, negedge CPN &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, negedge CPN &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, negedge CPN &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, negedge CPN &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, negedge CPN &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, negedge CPN &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNSND1 (SI, D, SE, CPN, SDN, Q, QN);
    input SI, D, SE, CPN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CPN_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_SE_SI_SDFCHK, CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_SI_SDFCHK, CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_nSI_SDFCHK, CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_SI_SDFCHK, CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SE_nSI_SDFCHK, CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_nSI_SDFCHK, CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_SI_SDFCHK, CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_nSI_SDFCHK, CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_SI_SDFCHK, nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_nSI_SDFCHK, nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_SI_SDFCHK, nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_nSI_SDFCHK, nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_SI_SDFCHK, nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_nSI_SDFCHK, nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_SI_SDFCHK, nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_nSI_SDFCHK, nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCPN, CPN);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CPN_D_SE_SI, CPN, D, SE, SI);
    and (CPN_D_nSE_SI, CPN, D, nSE, SI);
    and (CPN_D_nSE_nSI, CPN, D, nSE, nSI);
    and (CPN_nD_SE_SI, CPN, nD, SE, SI);
    and (CPN_D_SE_nSI, CPN, D, SE, nSI);
    and (CPN_nD_SE_nSI, CPN, nD, SE, nSI);
    and (CPN_nD_nSE_SI, CPN, nD, nSE, SI);
    and (CPN_nD_nSE_nSI, CPN, nD, nSE, nSI);
    and (nCPN_D_SE_SI, nCPN, D, SE, SI);
    and (nCPN_D_SE_nSI, nCPN, D, SE, nSI);
    and (nCPN_D_nSE_SI, nCPN, D, nSE, SI);
    and (nCPN_D_nSE_nSI, nCPN, D, nSE, nSI);
    and (nCPN_nD_SE_SI, nCPN, nD, SE, SI);
    and (nCPN_nD_SE_nSI, nCPN, nD, SE, nSI);
    and (nCPN_nD_nSE_SI, nCPN, nD, nSE, SI);
    and (nCPN_nD_nSE_nSI, nCPN, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, SDN_i, SE);
  `endif
  and  (D_check, SDN_i, SE_int_not);
  buf  (CPN_check, SDN_i);
  buf  (SE_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, negedge CPN &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, negedge CPN &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, negedge CPN &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, negedge CPN &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, negedge CPN &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, negedge CPN &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, negedge CPN &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, negedge CPN &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, negedge CPN &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, negedge CPN &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, negedge CPN &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, negedge CPN &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNSND2 (SI, D, SE, CPN, SDN, Q, QN);
    input SI, D, SE, CPN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CPN_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_SE_SI_SDFCHK, CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_SI_SDFCHK, CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_nSI_SDFCHK, CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_SI_SDFCHK, CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SE_nSI_SDFCHK, CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_nSI_SDFCHK, CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_SI_SDFCHK, CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_nSI_SDFCHK, CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_SI_SDFCHK, nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_nSI_SDFCHK, nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_SI_SDFCHK, nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_nSI_SDFCHK, nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_SI_SDFCHK, nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_nSI_SDFCHK, nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_SI_SDFCHK, nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_nSI_SDFCHK, nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCPN, CPN);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CPN_D_SE_SI, CPN, D, SE, SI);
    and (CPN_D_nSE_SI, CPN, D, nSE, SI);
    and (CPN_D_nSE_nSI, CPN, D, nSE, nSI);
    and (CPN_nD_SE_SI, CPN, nD, SE, SI);
    and (CPN_D_SE_nSI, CPN, D, SE, nSI);
    and (CPN_nD_SE_nSI, CPN, nD, SE, nSI);
    and (CPN_nD_nSE_SI, CPN, nD, nSE, SI);
    and (CPN_nD_nSE_nSI, CPN, nD, nSE, nSI);
    and (nCPN_D_SE_SI, nCPN, D, SE, SI);
    and (nCPN_D_SE_nSI, nCPN, D, SE, nSI);
    and (nCPN_D_nSE_SI, nCPN, D, nSE, SI);
    and (nCPN_D_nSE_nSI, nCPN, D, nSE, nSI);
    and (nCPN_nD_SE_SI, nCPN, nD, SE, SI);
    and (nCPN_nD_SE_nSI, nCPN, nD, SE, nSI);
    and (nCPN_nD_nSE_SI, nCPN, nD, nSE, SI);
    and (nCPN_nD_nSE_nSI, nCPN, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, SDN_i, SE);
  `endif
  and  (D_check, SDN_i, SE_int_not);
  buf  (CPN_check, SDN_i);
  buf  (SE_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, negedge CPN &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, negedge CPN &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, negedge CPN &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, negedge CPN &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, negedge CPN &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, negedge CPN &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, negedge CPN &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, negedge CPN &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, negedge CPN &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, negedge CPN &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, negedge CPN &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, negedge CPN &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNSND4 (SI, D, SE, CPN, SDN, Q, QN);
    input SI, D, SE, CPN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CPN_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_SE_SI_SDFCHK, CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_SI_SDFCHK, CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_nSI_SDFCHK, CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_SI_SDFCHK, CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SE_nSI_SDFCHK, CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_nSI_SDFCHK, CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_SI_SDFCHK, CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_nSI_SDFCHK, CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_SI_SDFCHK, nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_nSI_SDFCHK, nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_SI_SDFCHK, nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_nSI_SDFCHK, nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_SI_SDFCHK, nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_nSI_SDFCHK, nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_SI_SDFCHK, nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_nSI_SDFCHK, nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCPN, CPN);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CPN_D_SE_SI, CPN, D, SE, SI);
    and (CPN_D_nSE_SI, CPN, D, nSE, SI);
    and (CPN_D_nSE_nSI, CPN, D, nSE, nSI);
    and (CPN_nD_SE_SI, CPN, nD, SE, SI);
    and (CPN_D_SE_nSI, CPN, D, SE, nSI);
    and (CPN_nD_SE_nSI, CPN, nD, SE, nSI);
    and (CPN_nD_nSE_SI, CPN, nD, nSE, SI);
    and (CPN_nD_nSE_nSI, CPN, nD, nSE, nSI);
    and (nCPN_D_SE_SI, nCPN, D, SE, SI);
    and (nCPN_D_SE_nSI, nCPN, D, SE, nSI);
    and (nCPN_D_nSE_SI, nCPN, D, nSE, SI);
    and (nCPN_D_nSE_nSI, nCPN, D, nSE, nSI);
    and (nCPN_nD_SE_SI, nCPN, nD, SE, SI);
    and (nCPN_nD_SE_nSI, nCPN, nD, SE, nSI);
    and (nCPN_nD_nSE_SI, nCPN, nD, nSE, SI);
    and (nCPN_nD_nSE_nSI, nCPN, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, SDN_i, SE);
  `endif
  and  (D_check, SDN_i, SE_int_not);
  buf  (CPN_check, SDN_i);
  buf  (SE_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, negedge CPN &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, negedge CPN &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, negedge CPN &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, negedge CPN &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, negedge CPN &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, negedge CPN &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, negedge CPN &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, negedge CPN &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, negedge CPN &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, negedge CPN &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, negedge CPN &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, negedge CPN &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFQD0 (SI, D, SE, CP, Q);
    input SI, D, SE, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CP_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFQD1 (SI, D, SE, CP, Q);
    input SI, D, SE, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CP_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFQD2 (SI, D, SE, CP, Q);
    input SI, D, SE, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CP_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFQD4 (SI, D, SE, CP, Q);
    input SI, D, SE, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CP_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFQND0 (SI, D, SE, CP, QN);
    input SI, D, SE, CP;
    output QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (D_nSI, D, nSI);
    and (nD_SI, nD, SI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CP_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFQND1 (SI, D, SE, CP, QN);
    input SI, D, SE, CP;
    output QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (D_nSI, D, nSI);
    and (nD_SI, nD, SI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CP_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFQND2 (SI, D, SE, CP, QN);
    input SI, D, SE, CP;
    output QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (D_nSI, D, nSI);
    and (nD_SI, nD, SI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CP_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFQND4 (SI, D, SE, CP, QN);
    input SI, D, SE, CP;
    output QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (D_nSI, D, nSI);
    and (nD_SI, nD, SI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CP_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSND0 (SI, D, SE, CP, SDN, Q, QN);
    input SI, D, SE, CP, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, SDN_i, SE);
  `endif
  and  (D_check, SDN_i, SE_int_not);
  buf  (CP_check, SDN_i);
  buf  (SE_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSND1 (SI, D, SE, CP, SDN, Q, QN);
    input SI, D, SE, CP, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, SDN_i, SE);
  `endif
  and  (D_check, SDN_i, SE_int_not);
  buf  (CP_check, SDN_i);
  buf  (SE_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSND2 (SI, D, SE, CP, SDN, Q, QN);
    input SI, D, SE, CP, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, SDN_i, SE);
  `endif
  and  (D_check, SDN_i, SE_int_not);
  buf  (CP_check, SDN_i);
  buf  (SE_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSND4 (SI, D, SE, CP, SDN, Q, QN);
    input SI, D, SE, CP, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, SDN_i, SE);
  `endif
  and  (D_check, SDN_i, SE_int_not);
  buf  (CP_check, SDN_i);
  buf  (SE_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSNQD0 (SI, D, SE, CP, SDN, Q);
    input SI, D, SE, CP, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, SDN_i, SE);
  `endif
  and  (D_check, SDN_i, SE_int_not);
  buf  (CP_check, SDN_i);
  buf  (SE_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSNQD1 (SI, D, SE, CP, SDN, Q);
    input SI, D, SE, CP, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, SDN_i, SE);
  `endif
  and  (D_check, SDN_i, SE_int_not);
  buf  (CP_check, SDN_i);
  buf  (SE_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSNQD2 (SI, D, SE, CP, SDN, Q);
    input SI, D, SE, CP, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, SDN_i, SE);
  `endif
  and  (D_check, SDN_i, SE_int_not);
  buf  (CP_check, SDN_i);
  buf  (SE_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSNQD4 (SI, D, SE, CP, SDN, Q);
    input SI, D, SE, CP, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, SDN_i, SE);
  `endif
  and  (D_check, SDN_i, SE_int_not);
  buf  (CP_check, SDN_i);
  buf  (SE_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFXD0 (DA, DB, SA, SI, SE, CP, Q, QN);
    input DA, DB, SA, SI, SE, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire DA_d, DB_d, SA_d, SI_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB_d, DA_d, SA_d);
        tsmc_mux (D_i, D, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB, DA, SA);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (DA_DB_SA_SE_SI_SDFCHK, DA_DB_SA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSE_SI_SDFCHK, DA_DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSE_nSI_SDFCHK, DA_DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_SI_SDFCHK, DA_DB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSE_SI_SDFCHK, DA_DB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSE_nSI_SDFCHK, DA_DB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_SI_SDFCHK, DA_nDB_SA_SE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSE_SI_SDFCHK, DA_nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSE_nSI_SDFCHK, DA_nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_SI_SDFCHK, DA_nDB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_SI_SDFCHK, nDA_DB_SA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_SI_SDFCHK, nDA_DB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSE_SI_SDFCHK, nDA_DB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSE_nSI_SDFCHK, nDA_DB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_SI_SDFCHK, nDA_nDB_SA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_SI_SDFCHK, nDA_nDB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_SE_nSI_SDFCHK, DA_DB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_nSI_SDFCHK, DA_DB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_nSI_SDFCHK, DA_nDB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_nSI_SDFCHK, DA_nDB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_nSE_SI_SDFCHK, DA_nDB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_nSE_nSI_SDFCHK, DA_nDB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_nSI_SDFCHK, nDA_DB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_nSE_SI_SDFCHK, nDA_DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_nSE_nSI_SDFCHK, nDA_DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_nSI_SDFCHK, nDA_DB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_nSI_SDFCHK, nDA_nDB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_nSE_SI_SDFCHK, nDA_nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_nSE_nSI_SDFCHK, nDA_nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_nSI_SDFCHK, nDA_nDB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_nSE_SI_SDFCHK, nDA_nDB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_nSE_nSI_SDFCHK, nDA_nDB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DB_SA_nSE_SI_SDFCHK, DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DB_SA_nSE_nSI_SDFCHK, DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDB_SA_nSE_SI_SDFCHK, nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDB_SA_nSE_nSI_SDFCHK, nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nSA_nSE_SI_SDFCHK, DA_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nSA_nSE_nSI_SDFCHK, DA_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nSA_nSE_SI_SDFCHK, nDA_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nSA_nSE_nSI_SDFCHK, nDA_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSE_SI_SDFCHK, DA_nDB_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_nSE_nSI_SDFCHK, DA_nDB_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSE_SI_SDFCHK, nDA_DB_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSE_nSI_SDFCHK, nDA_DB_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SI_SDFCHK, DA_nDB_nSA_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SI_SDFCHK, nDA_DB_SA_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SI_SDFCHK, nDA_nDB_SA_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SI_SDFCHK, nDA_nDB_nSA_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSI_SDFCHK, DA_DB_SA_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSI_SDFCHK, DA_DB_nSA_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSI_SDFCHK, DA_nDB_SA_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSI_SDFCHK, nDA_DB_nSA_nSI, 1'b1);
    tsmc_xbuf (DA_DB_SA_SE_SDFCHK, DA_DB_SA_SE, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_SDFCHK, DA_DB_nSA_SE, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_SDFCHK, DA_nDB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_SDFCHK, nDA_DB_nSA_SE, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_SDFCHK, DA_nDB_nSA_SE, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_SDFCHK, nDA_DB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_SDFCHK, nDA_nDB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_SDFCHK, nDA_nDB_nSA_SE, 1'b1);
  `endif

    not (nDA, DA);
    not (nDB, DB);
    not (nSA, SA);
    not (nSI, SI);
    not (nSE, SE);
    and (DA_DB_SA_SE_SI, DA, DB, SA, SE, SI);
    and (DA_DB_SA_nSE_SI, DA, DB, SA, nSE, SI);
    and (DA_DB_SA_nSE_nSI, DA, DB, SA, nSE, nSI);
    and (DA_DB_nSA_SE_SI, DA, DB, nSA, SE, SI);
    and (DA_DB_nSA_nSE_SI, DA, DB, nSA, nSE, SI);
    and (DA_DB_nSA_nSE_nSI, DA, DB, nSA, nSE, nSI);
    and (DA_nDB_SA_SE_SI, DA, nDB, SA, SE, SI);
    and (DA_nDB_SA_nSE_SI, DA, nDB, SA, nSE, SI);
    and (DA_nDB_SA_nSE_nSI, DA, nDB, SA, nSE, nSI);
    and (DA_nDB_nSA_SE_SI, DA, nDB, nSA, SE, SI);
    and (nDA_DB_SA_SE_SI, nDA, DB, SA, SE, SI);
    and (nDA_DB_nSA_SE_SI, nDA, DB, nSA, SE, SI);
    and (nDA_DB_nSA_nSE_SI, nDA, DB, nSA, nSE, SI);
    and (nDA_DB_nSA_nSE_nSI, nDA, DB, nSA, nSE, nSI);
    and (nDA_nDB_SA_SE_SI, nDA, nDB, SA, SE, SI);
    and (nDA_nDB_nSA_SE_SI, nDA, nDB, nSA, SE, SI);
    and (DA_DB_SA_SE_nSI, DA, DB, SA, SE, nSI);
    and (DA_DB_nSA_SE_nSI, DA, DB, nSA, SE, nSI);
    and (DA_nDB_SA_SE_nSI, DA, nDB, SA, SE, nSI);
    and (DA_nDB_nSA_SE_nSI, DA, nDB, nSA, SE, nSI);
    and (DA_nDB_nSA_nSE_SI, DA, nDB, nSA, nSE, SI);
    and (DA_nDB_nSA_nSE_nSI, DA, nDB, nSA, nSE, nSI);
    and (nDA_DB_SA_SE_nSI, nDA, DB, SA, SE, nSI);
    and (nDA_DB_SA_nSE_SI, nDA, DB, SA, nSE, SI);
    and (nDA_DB_SA_nSE_nSI, nDA, DB, SA, nSE, nSI);
    and (nDA_DB_nSA_SE_nSI, nDA, DB, nSA, SE, nSI);
    and (nDA_nDB_SA_SE_nSI, nDA, nDB, SA, SE, nSI);
    and (nDA_nDB_SA_nSE_SI, nDA, nDB, SA, nSE, SI);
    and (nDA_nDB_SA_nSE_nSI, nDA, nDB, SA, nSE, nSI);
    and (nDA_nDB_nSA_SE_nSI, nDA, nDB, nSA, SE, nSI);
    and (nDA_nDB_nSA_nSE_SI, nDA, nDB, nSA, nSE, SI);
    and (nDA_nDB_nSA_nSE_nSI, nDA, nDB, nSA, nSE, nSI);
    and (DB_SA_nSE_SI, DB, SA, nSE, SI);
    and (DB_SA_nSE_nSI, DB, SA, nSE, nSI);
    and (nDB_SA_nSE_SI, nDB, SA, nSE, SI);
    and (nDB_SA_nSE_nSI, nDB, SA, nSE, nSI);
    and (DA_nSA_nSE_SI, DA, nSA, nSE, SI);
    and (DA_nSA_nSE_nSI, DA, nSA, nSE, nSI);
    and (nDA_nSA_nSE_SI, nDA, nSA, nSE, SI);
    and (nDA_nSA_nSE_nSI, nDA, nSA, nSE, nSI);
    and (DA_nDB_nSE_SI, DA, nDB, nSE, SI);
    and (DA_nDB_nSE_nSI, DA, nDB, nSE, nSI);
    and (nDA_DB_nSE_SI, nDA, DB, nSE, SI);
    and (nDA_DB_nSE_nSI, nDA, DB, nSE, nSI);
    and (DA_nDB_nSA_SI, DA, nDB, nSA, SI);
    and (nDA_DB_SA_SI, nDA, DB, SA, SI);
    and (nDA_nDB_SA_SI, nDA, nDB, SA, SI);
    and (nDA_nDB_nSA_SI, nDA, nDB, nSA, SI);
    and (DA_DB_SA_nSI, DA, DB, SA, nSI);
    and (DA_DB_nSA_nSI, DA, DB, nSA, nSI);
    and (DA_nDB_SA_nSI, DA, nDB, SA, nSI);
    and (nDA_DB_nSA_nSI, nDA, DB, nSA, nSI);
    and (DA_DB_SA_SE, DA, DB, SA, SE);
    and (DA_DB_nSA_SE, DA, DB, nSA, SE);
    and (DA_nDB_SA_SE, DA, nDB, SA, SE);
    and (nDA_DB_nSA_SE, nDA, DB, nSA, SE);
    and (DA_nDB_nSA_SE, DA, nDB, nSA, SE);
    and (nDA_DB_SA_SE, nDA, DB, SA, SE);
    and (nDA_nDB_SA_SE, nDA, nDB, SA, SE);
    and (nDA_nDB_nSA_SE, nDA, nDB, nSA, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SA_int_not, SA_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (DA_check, SA_d, SE_int_not);
  `else
    not  (SA_int_not, SA);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (DA_check, SA, SE_int_not);
  `endif
  buf  (SA_check, SE_int_not);
  and  (DB_check, SA_int_not, SE_int_not);
  or   (CP_check, SI_check, DA_check, SA_check, DB_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    $width (posedge CP &&& DA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFXD1 (DA, DB, SA, SI, SE, CP, Q, QN);
    input DA, DB, SA, SI, SE, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire DA_d, DB_d, SA_d, SI_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB_d, DA_d, SA_d);
        tsmc_mux (D_i, D, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB, DA, SA);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (DA_DB_SA_SE_SI_SDFCHK, DA_DB_SA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSE_SI_SDFCHK, DA_DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSE_nSI_SDFCHK, DA_DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_SI_SDFCHK, DA_DB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSE_SI_SDFCHK, DA_DB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSE_nSI_SDFCHK, DA_DB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_SI_SDFCHK, DA_nDB_SA_SE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSE_SI_SDFCHK, DA_nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSE_nSI_SDFCHK, DA_nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_SI_SDFCHK, DA_nDB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_SI_SDFCHK, nDA_DB_SA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_SI_SDFCHK, nDA_DB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSE_SI_SDFCHK, nDA_DB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSE_nSI_SDFCHK, nDA_DB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_SI_SDFCHK, nDA_nDB_SA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_SI_SDFCHK, nDA_nDB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_SE_nSI_SDFCHK, DA_DB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_nSI_SDFCHK, DA_DB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_nSI_SDFCHK, DA_nDB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_nSI_SDFCHK, DA_nDB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_nSE_SI_SDFCHK, DA_nDB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_nSE_nSI_SDFCHK, DA_nDB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_nSI_SDFCHK, nDA_DB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_nSE_SI_SDFCHK, nDA_DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_nSE_nSI_SDFCHK, nDA_DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_nSI_SDFCHK, nDA_DB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_nSI_SDFCHK, nDA_nDB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_nSE_SI_SDFCHK, nDA_nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_nSE_nSI_SDFCHK, nDA_nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_nSI_SDFCHK, nDA_nDB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_nSE_SI_SDFCHK, nDA_nDB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_nSE_nSI_SDFCHK, nDA_nDB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DB_SA_nSE_SI_SDFCHK, DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DB_SA_nSE_nSI_SDFCHK, DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDB_SA_nSE_SI_SDFCHK, nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDB_SA_nSE_nSI_SDFCHK, nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nSA_nSE_SI_SDFCHK, DA_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nSA_nSE_nSI_SDFCHK, DA_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nSA_nSE_SI_SDFCHK, nDA_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nSA_nSE_nSI_SDFCHK, nDA_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSE_SI_SDFCHK, DA_nDB_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_nSE_nSI_SDFCHK, DA_nDB_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSE_SI_SDFCHK, nDA_DB_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSE_nSI_SDFCHK, nDA_DB_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SI_SDFCHK, DA_nDB_nSA_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SI_SDFCHK, nDA_DB_SA_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SI_SDFCHK, nDA_nDB_SA_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SI_SDFCHK, nDA_nDB_nSA_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSI_SDFCHK, DA_DB_SA_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSI_SDFCHK, DA_DB_nSA_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSI_SDFCHK, DA_nDB_SA_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSI_SDFCHK, nDA_DB_nSA_nSI, 1'b1);
    tsmc_xbuf (DA_DB_SA_SE_SDFCHK, DA_DB_SA_SE, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_SDFCHK, DA_DB_nSA_SE, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_SDFCHK, DA_nDB_SA_SE, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_SDFCHK, DA_nDB_nSA_SE, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_SDFCHK, nDA_DB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_SDFCHK, nDA_DB_nSA_SE, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_SDFCHK, nDA_nDB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_SDFCHK, nDA_nDB_nSA_SE, 1'b1);
  `endif

    not (nDA, DA);
    not (nDB, DB);
    not (nSA, SA);
    not (nSI, SI);
    not (nSE, SE);
    and (DA_DB_SA_SE_SI, DA, DB, SA, SE, SI);
    and (DA_DB_SA_nSE_SI, DA, DB, SA, nSE, SI);
    and (DA_DB_SA_nSE_nSI, DA, DB, SA, nSE, nSI);
    and (DA_DB_nSA_SE_SI, DA, DB, nSA, SE, SI);
    and (DA_DB_nSA_nSE_SI, DA, DB, nSA, nSE, SI);
    and (DA_DB_nSA_nSE_nSI, DA, DB, nSA, nSE, nSI);
    and (DA_nDB_SA_SE_SI, DA, nDB, SA, SE, SI);
    and (DA_nDB_SA_nSE_SI, DA, nDB, SA, nSE, SI);
    and (DA_nDB_SA_nSE_nSI, DA, nDB, SA, nSE, nSI);
    and (DA_nDB_nSA_SE_SI, DA, nDB, nSA, SE, SI);
    and (nDA_DB_SA_SE_SI, nDA, DB, SA, SE, SI);
    and (nDA_DB_nSA_SE_SI, nDA, DB, nSA, SE, SI);
    and (nDA_DB_nSA_nSE_SI, nDA, DB, nSA, nSE, SI);
    and (nDA_DB_nSA_nSE_nSI, nDA, DB, nSA, nSE, nSI);
    and (nDA_nDB_SA_SE_SI, nDA, nDB, SA, SE, SI);
    and (nDA_nDB_nSA_SE_SI, nDA, nDB, nSA, SE, SI);
    and (DA_DB_SA_SE_nSI, DA, DB, SA, SE, nSI);
    and (DA_DB_nSA_SE_nSI, DA, DB, nSA, SE, nSI);
    and (DA_nDB_SA_SE_nSI, DA, nDB, SA, SE, nSI);
    and (DA_nDB_nSA_SE_nSI, DA, nDB, nSA, SE, nSI);
    and (DA_nDB_nSA_nSE_SI, DA, nDB, nSA, nSE, SI);
    and (DA_nDB_nSA_nSE_nSI, DA, nDB, nSA, nSE, nSI);
    and (nDA_DB_SA_SE_nSI, nDA, DB, SA, SE, nSI);
    and (nDA_DB_SA_nSE_SI, nDA, DB, SA, nSE, SI);
    and (nDA_DB_SA_nSE_nSI, nDA, DB, SA, nSE, nSI);
    and (nDA_DB_nSA_SE_nSI, nDA, DB, nSA, SE, nSI);
    and (nDA_nDB_SA_SE_nSI, nDA, nDB, SA, SE, nSI);
    and (nDA_nDB_SA_nSE_SI, nDA, nDB, SA, nSE, SI);
    and (nDA_nDB_SA_nSE_nSI, nDA, nDB, SA, nSE, nSI);
    and (nDA_nDB_nSA_SE_nSI, nDA, nDB, nSA, SE, nSI);
    and (nDA_nDB_nSA_nSE_SI, nDA, nDB, nSA, nSE, SI);
    and (nDA_nDB_nSA_nSE_nSI, nDA, nDB, nSA, nSE, nSI);
    and (DB_SA_nSE_SI, DB, SA, nSE, SI);
    and (DB_SA_nSE_nSI, DB, SA, nSE, nSI);
    and (nDB_SA_nSE_SI, nDB, SA, nSE, SI);
    and (nDB_SA_nSE_nSI, nDB, SA, nSE, nSI);
    and (DA_nSA_nSE_SI, DA, nSA, nSE, SI);
    and (DA_nSA_nSE_nSI, DA, nSA, nSE, nSI);
    and (nDA_nSA_nSE_SI, nDA, nSA, nSE, SI);
    and (nDA_nSA_nSE_nSI, nDA, nSA, nSE, nSI);
    and (DA_nDB_nSE_SI, DA, nDB, nSE, SI);
    and (DA_nDB_nSE_nSI, DA, nDB, nSE, nSI);
    and (nDA_DB_nSE_SI, nDA, DB, nSE, SI);
    and (nDA_DB_nSE_nSI, nDA, DB, nSE, nSI);
    and (DA_nDB_nSA_SI, DA, nDB, nSA, SI);
    and (nDA_DB_SA_SI, nDA, DB, SA, SI);
    and (nDA_nDB_SA_SI, nDA, nDB, SA, SI);
    and (nDA_nDB_nSA_SI, nDA, nDB, nSA, SI);
    and (DA_DB_SA_nSI, DA, DB, SA, nSI);
    and (DA_DB_nSA_nSI, DA, DB, nSA, nSI);
    and (DA_nDB_SA_nSI, DA, nDB, SA, nSI);
    and (nDA_DB_nSA_nSI, nDA, DB, nSA, nSI);
    and (DA_DB_SA_SE, DA, DB, SA, SE);
    and (DA_DB_nSA_SE, DA, DB, nSA, SE);
    and (DA_nDB_SA_SE, DA, nDB, SA, SE);
    and (DA_nDB_nSA_SE, DA, nDB, nSA, SE);
    and (nDA_DB_SA_SE, nDA, DB, SA, SE);
    and (nDA_DB_nSA_SE, nDA, DB, nSA, SE);
    and (nDA_nDB_SA_SE, nDA, nDB, SA, SE);
    and (nDA_nDB_nSA_SE, nDA, nDB, nSA, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SA_int_not, SA_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (DA_check, SA_d, SE_int_not);
  `else
    not  (SA_int_not, SA);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (DA_check, SA, SE_int_not);
  `endif
  buf  (SA_check, SE_int_not);
  and  (DB_check, SA_int_not, SE_int_not);
  or   (CP_check, SI_check, DA_check, SA_check, DB_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    $width (posedge CP &&& DA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFXD2 (DA, DB, SA, SI, SE, CP, Q, QN);
    input DA, DB, SA, SI, SE, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire DA_d, DB_d, SA_d, SI_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB_d, DA_d, SA_d);
        tsmc_mux (D_i, D, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB, DA, SA);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (DA_DB_SA_SE_SI_SDFCHK, DA_DB_SA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSE_SI_SDFCHK, DA_DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSE_nSI_SDFCHK, DA_DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_SI_SDFCHK, DA_DB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSE_SI_SDFCHK, DA_DB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSE_nSI_SDFCHK, DA_DB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_SI_SDFCHK, DA_nDB_SA_SE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSE_SI_SDFCHK, DA_nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSE_nSI_SDFCHK, DA_nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_SI_SDFCHK, DA_nDB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_SI_SDFCHK, nDA_DB_SA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_SI_SDFCHK, nDA_DB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSE_SI_SDFCHK, nDA_DB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSE_nSI_SDFCHK, nDA_DB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_SI_SDFCHK, nDA_nDB_SA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_SI_SDFCHK, nDA_nDB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_SE_nSI_SDFCHK, DA_DB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_nSI_SDFCHK, DA_DB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_nSI_SDFCHK, DA_nDB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_nSI_SDFCHK, DA_nDB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_nSE_SI_SDFCHK, DA_nDB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_nSE_nSI_SDFCHK, DA_nDB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_nSI_SDFCHK, nDA_DB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_nSE_SI_SDFCHK, nDA_DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_nSE_nSI_SDFCHK, nDA_DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_nSI_SDFCHK, nDA_DB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_nSI_SDFCHK, nDA_nDB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_nSE_SI_SDFCHK, nDA_nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_nSE_nSI_SDFCHK, nDA_nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_nSI_SDFCHK, nDA_nDB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_nSE_SI_SDFCHK, nDA_nDB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_nSE_nSI_SDFCHK, nDA_nDB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DB_SA_nSE_SI_SDFCHK, DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DB_SA_nSE_nSI_SDFCHK, DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDB_SA_nSE_SI_SDFCHK, nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDB_SA_nSE_nSI_SDFCHK, nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nSA_nSE_SI_SDFCHK, DA_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nSA_nSE_nSI_SDFCHK, DA_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nSA_nSE_SI_SDFCHK, nDA_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nSA_nSE_nSI_SDFCHK, nDA_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSE_SI_SDFCHK, DA_nDB_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_nSE_nSI_SDFCHK, DA_nDB_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSE_SI_SDFCHK, nDA_DB_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSE_nSI_SDFCHK, nDA_DB_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SI_SDFCHK, DA_nDB_nSA_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SI_SDFCHK, nDA_DB_SA_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SI_SDFCHK, nDA_nDB_SA_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SI_SDFCHK, nDA_nDB_nSA_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSI_SDFCHK, DA_DB_SA_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSI_SDFCHK, DA_DB_nSA_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSI_SDFCHK, DA_nDB_SA_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSI_SDFCHK, nDA_DB_nSA_nSI, 1'b1);
    tsmc_xbuf (DA_DB_SA_SE_SDFCHK, DA_DB_SA_SE, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_SDFCHK, DA_DB_nSA_SE, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_SDFCHK, DA_nDB_SA_SE, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_SDFCHK, DA_nDB_nSA_SE, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_SDFCHK, nDA_DB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_SDFCHK, nDA_DB_nSA_SE, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_SDFCHK, nDA_nDB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_SDFCHK, nDA_nDB_nSA_SE, 1'b1);
  `endif

    not (nDA, DA);
    not (nDB, DB);
    not (nSA, SA);
    not (nSI, SI);
    not (nSE, SE);
    and (DA_DB_SA_SE_SI, DA, DB, SA, SE, SI);
    and (DA_DB_SA_nSE_SI, DA, DB, SA, nSE, SI);
    and (DA_DB_SA_nSE_nSI, DA, DB, SA, nSE, nSI);
    and (DA_DB_nSA_SE_SI, DA, DB, nSA, SE, SI);
    and (DA_DB_nSA_nSE_SI, DA, DB, nSA, nSE, SI);
    and (DA_DB_nSA_nSE_nSI, DA, DB, nSA, nSE, nSI);
    and (DA_nDB_SA_SE_SI, DA, nDB, SA, SE, SI);
    and (DA_nDB_SA_nSE_SI, DA, nDB, SA, nSE, SI);
    and (DA_nDB_SA_nSE_nSI, DA, nDB, SA, nSE, nSI);
    and (DA_nDB_nSA_SE_SI, DA, nDB, nSA, SE, SI);
    and (nDA_DB_SA_SE_SI, nDA, DB, SA, SE, SI);
    and (nDA_DB_nSA_SE_SI, nDA, DB, nSA, SE, SI);
    and (nDA_DB_nSA_nSE_SI, nDA, DB, nSA, nSE, SI);
    and (nDA_DB_nSA_nSE_nSI, nDA, DB, nSA, nSE, nSI);
    and (nDA_nDB_SA_SE_SI, nDA, nDB, SA, SE, SI);
    and (nDA_nDB_nSA_SE_SI, nDA, nDB, nSA, SE, SI);
    and (DA_DB_SA_SE_nSI, DA, DB, SA, SE, nSI);
    and (DA_DB_nSA_SE_nSI, DA, DB, nSA, SE, nSI);
    and (DA_nDB_SA_SE_nSI, DA, nDB, SA, SE, nSI);
    and (DA_nDB_nSA_SE_nSI, DA, nDB, nSA, SE, nSI);
    and (DA_nDB_nSA_nSE_SI, DA, nDB, nSA, nSE, SI);
    and (DA_nDB_nSA_nSE_nSI, DA, nDB, nSA, nSE, nSI);
    and (nDA_DB_SA_SE_nSI, nDA, DB, SA, SE, nSI);
    and (nDA_DB_SA_nSE_SI, nDA, DB, SA, nSE, SI);
    and (nDA_DB_SA_nSE_nSI, nDA, DB, SA, nSE, nSI);
    and (nDA_DB_nSA_SE_nSI, nDA, DB, nSA, SE, nSI);
    and (nDA_nDB_SA_SE_nSI, nDA, nDB, SA, SE, nSI);
    and (nDA_nDB_SA_nSE_SI, nDA, nDB, SA, nSE, SI);
    and (nDA_nDB_SA_nSE_nSI, nDA, nDB, SA, nSE, nSI);
    and (nDA_nDB_nSA_SE_nSI, nDA, nDB, nSA, SE, nSI);
    and (nDA_nDB_nSA_nSE_SI, nDA, nDB, nSA, nSE, SI);
    and (nDA_nDB_nSA_nSE_nSI, nDA, nDB, nSA, nSE, nSI);
    and (DB_SA_nSE_SI, DB, SA, nSE, SI);
    and (DB_SA_nSE_nSI, DB, SA, nSE, nSI);
    and (nDB_SA_nSE_SI, nDB, SA, nSE, SI);
    and (nDB_SA_nSE_nSI, nDB, SA, nSE, nSI);
    and (DA_nSA_nSE_SI, DA, nSA, nSE, SI);
    and (DA_nSA_nSE_nSI, DA, nSA, nSE, nSI);
    and (nDA_nSA_nSE_SI, nDA, nSA, nSE, SI);
    and (nDA_nSA_nSE_nSI, nDA, nSA, nSE, nSI);
    and (DA_nDB_nSE_SI, DA, nDB, nSE, SI);
    and (DA_nDB_nSE_nSI, DA, nDB, nSE, nSI);
    and (nDA_DB_nSE_SI, nDA, DB, nSE, SI);
    and (nDA_DB_nSE_nSI, nDA, DB, nSE, nSI);
    and (DA_nDB_nSA_SI, DA, nDB, nSA, SI);
    and (nDA_DB_SA_SI, nDA, DB, SA, SI);
    and (nDA_nDB_SA_SI, nDA, nDB, SA, SI);
    and (nDA_nDB_nSA_SI, nDA, nDB, nSA, SI);
    and (DA_DB_SA_nSI, DA, DB, SA, nSI);
    and (DA_DB_nSA_nSI, DA, DB, nSA, nSI);
    and (DA_nDB_SA_nSI, DA, nDB, SA, nSI);
    and (nDA_DB_nSA_nSI, nDA, DB, nSA, nSI);
    and (DA_DB_SA_SE, DA, DB, SA, SE);
    and (DA_DB_nSA_SE, DA, DB, nSA, SE);
    and (DA_nDB_SA_SE, DA, nDB, SA, SE);
    and (DA_nDB_nSA_SE, DA, nDB, nSA, SE);
    and (nDA_DB_SA_SE, nDA, DB, SA, SE);
    and (nDA_DB_nSA_SE, nDA, DB, nSA, SE);
    and (nDA_nDB_SA_SE, nDA, nDB, SA, SE);
    and (nDA_nDB_nSA_SE, nDA, nDB, nSA, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SA_int_not, SA_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (DA_check, SA_d, SE_int_not);
  `else
    not  (SA_int_not, SA);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (DA_check, SA, SE_int_not);
  `endif
  buf  (SA_check, SE_int_not);
  and  (DB_check, SA_int_not, SE_int_not);
  or   (CP_check, SI_check, DA_check, SA_check, DB_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    $width (posedge CP &&& DA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFXD4 (DA, DB, SA, SI, SE, CP, Q, QN);
    input DA, DB, SA, SI, SE, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire DA_d, DB_d, SA_d, SI_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB_d, DA_d, SA_d);
        tsmc_mux (D_i, D, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB, DA, SA);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (DA_DB_SA_SE_SI_SDFCHK, DA_DB_SA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSE_SI_SDFCHK, DA_DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSE_nSI_SDFCHK, DA_DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_SI_SDFCHK, DA_DB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSE_SI_SDFCHK, DA_DB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSE_nSI_SDFCHK, DA_DB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_SI_SDFCHK, DA_nDB_SA_SE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSE_SI_SDFCHK, DA_nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSE_nSI_SDFCHK, DA_nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_SI_SDFCHK, DA_nDB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_SI_SDFCHK, nDA_DB_SA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_SI_SDFCHK, nDA_DB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSE_SI_SDFCHK, nDA_DB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSE_nSI_SDFCHK, nDA_DB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_SI_SDFCHK, nDA_nDB_SA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_SI_SDFCHK, nDA_nDB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_SE_nSI_SDFCHK, DA_DB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_nSI_SDFCHK, DA_DB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_nSI_SDFCHK, DA_nDB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_nSI_SDFCHK, DA_nDB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_nSE_SI_SDFCHK, DA_nDB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_nSE_nSI_SDFCHK, DA_nDB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_nSI_SDFCHK, nDA_DB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_nSE_SI_SDFCHK, nDA_DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_nSE_nSI_SDFCHK, nDA_DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_nSI_SDFCHK, nDA_DB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_nSI_SDFCHK, nDA_nDB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_nSE_SI_SDFCHK, nDA_nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_nSE_nSI_SDFCHK, nDA_nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_nSI_SDFCHK, nDA_nDB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_nSE_SI_SDFCHK, nDA_nDB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_nSE_nSI_SDFCHK, nDA_nDB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DB_SA_nSE_SI_SDFCHK, DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DB_SA_nSE_nSI_SDFCHK, DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDB_SA_nSE_SI_SDFCHK, nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDB_SA_nSE_nSI_SDFCHK, nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nSA_nSE_SI_SDFCHK, DA_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nSA_nSE_nSI_SDFCHK, DA_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nSA_nSE_SI_SDFCHK, nDA_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nSA_nSE_nSI_SDFCHK, nDA_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSE_SI_SDFCHK, DA_nDB_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_nSE_nSI_SDFCHK, DA_nDB_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSE_SI_SDFCHK, nDA_DB_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSE_nSI_SDFCHK, nDA_DB_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SI_SDFCHK, DA_nDB_nSA_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SI_SDFCHK, nDA_DB_SA_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SI_SDFCHK, nDA_nDB_SA_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SI_SDFCHK, nDA_nDB_nSA_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSI_SDFCHK, DA_DB_SA_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSI_SDFCHK, DA_DB_nSA_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSI_SDFCHK, DA_nDB_SA_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSI_SDFCHK, nDA_DB_nSA_nSI, 1'b1);
    tsmc_xbuf (DA_DB_SA_SE_SDFCHK, DA_DB_SA_SE, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_SDFCHK, DA_DB_nSA_SE, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_SDFCHK, DA_nDB_SA_SE, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_SDFCHK, DA_nDB_nSA_SE, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_SDFCHK, nDA_DB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_SDFCHK, nDA_DB_nSA_SE, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_SDFCHK, nDA_nDB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_SDFCHK, nDA_nDB_nSA_SE, 1'b1);
  `endif

    not (nDA, DA);
    not (nDB, DB);
    not (nSA, SA);
    not (nSI, SI);
    not (nSE, SE);
    and (DA_DB_SA_SE_SI, DA, DB, SA, SE, SI);
    and (DA_DB_SA_nSE_SI, DA, DB, SA, nSE, SI);
    and (DA_DB_SA_nSE_nSI, DA, DB, SA, nSE, nSI);
    and (DA_DB_nSA_SE_SI, DA, DB, nSA, SE, SI);
    and (DA_DB_nSA_nSE_SI, DA, DB, nSA, nSE, SI);
    and (DA_DB_nSA_nSE_nSI, DA, DB, nSA, nSE, nSI);
    and (DA_nDB_SA_SE_SI, DA, nDB, SA, SE, SI);
    and (DA_nDB_SA_nSE_SI, DA, nDB, SA, nSE, SI);
    and (DA_nDB_SA_nSE_nSI, DA, nDB, SA, nSE, nSI);
    and (DA_nDB_nSA_SE_SI, DA, nDB, nSA, SE, SI);
    and (nDA_DB_SA_SE_SI, nDA, DB, SA, SE, SI);
    and (nDA_DB_nSA_SE_SI, nDA, DB, nSA, SE, SI);
    and (nDA_DB_nSA_nSE_SI, nDA, DB, nSA, nSE, SI);
    and (nDA_DB_nSA_nSE_nSI, nDA, DB, nSA, nSE, nSI);
    and (nDA_nDB_SA_SE_SI, nDA, nDB, SA, SE, SI);
    and (nDA_nDB_nSA_SE_SI, nDA, nDB, nSA, SE, SI);
    and (DA_DB_SA_SE_nSI, DA, DB, SA, SE, nSI);
    and (DA_DB_nSA_SE_nSI, DA, DB, nSA, SE, nSI);
    and (DA_nDB_SA_SE_nSI, DA, nDB, SA, SE, nSI);
    and (DA_nDB_nSA_SE_nSI, DA, nDB, nSA, SE, nSI);
    and (DA_nDB_nSA_nSE_SI, DA, nDB, nSA, nSE, SI);
    and (DA_nDB_nSA_nSE_nSI, DA, nDB, nSA, nSE, nSI);
    and (nDA_DB_SA_SE_nSI, nDA, DB, SA, SE, nSI);
    and (nDA_DB_SA_nSE_SI, nDA, DB, SA, nSE, SI);
    and (nDA_DB_SA_nSE_nSI, nDA, DB, SA, nSE, nSI);
    and (nDA_DB_nSA_SE_nSI, nDA, DB, nSA, SE, nSI);
    and (nDA_nDB_SA_SE_nSI, nDA, nDB, SA, SE, nSI);
    and (nDA_nDB_SA_nSE_SI, nDA, nDB, SA, nSE, SI);
    and (nDA_nDB_SA_nSE_nSI, nDA, nDB, SA, nSE, nSI);
    and (nDA_nDB_nSA_SE_nSI, nDA, nDB, nSA, SE, nSI);
    and (nDA_nDB_nSA_nSE_SI, nDA, nDB, nSA, nSE, SI);
    and (nDA_nDB_nSA_nSE_nSI, nDA, nDB, nSA, nSE, nSI);
    and (DB_SA_nSE_SI, DB, SA, nSE, SI);
    and (DB_SA_nSE_nSI, DB, SA, nSE, nSI);
    and (nDB_SA_nSE_SI, nDB, SA, nSE, SI);
    and (nDB_SA_nSE_nSI, nDB, SA, nSE, nSI);
    and (DA_nSA_nSE_SI, DA, nSA, nSE, SI);
    and (DA_nSA_nSE_nSI, DA, nSA, nSE, nSI);
    and (nDA_nSA_nSE_SI, nDA, nSA, nSE, SI);
    and (nDA_nSA_nSE_nSI, nDA, nSA, nSE, nSI);
    and (DA_nDB_nSE_SI, DA, nDB, nSE, SI);
    and (DA_nDB_nSE_nSI, DA, nDB, nSE, nSI);
    and (nDA_DB_nSE_SI, nDA, DB, nSE, SI);
    and (nDA_DB_nSE_nSI, nDA, DB, nSE, nSI);
    and (DA_nDB_nSA_SI, DA, nDB, nSA, SI);
    and (nDA_DB_SA_SI, nDA, DB, SA, SI);
    and (nDA_nDB_SA_SI, nDA, nDB, SA, SI);
    and (nDA_nDB_nSA_SI, nDA, nDB, nSA, SI);
    and (DA_DB_SA_nSI, DA, DB, SA, nSI);
    and (DA_DB_nSA_nSI, DA, DB, nSA, nSI);
    and (DA_nDB_SA_nSI, DA, nDB, SA, nSI);
    and (nDA_DB_nSA_nSI, nDA, DB, nSA, nSI);
    and (DA_DB_SA_SE, DA, DB, SA, SE);
    and (DA_DB_nSA_SE, DA, DB, nSA, SE);
    and (DA_nDB_SA_SE, DA, nDB, SA, SE);
    and (DA_nDB_nSA_SE, DA, nDB, nSA, SE);
    and (nDA_DB_SA_SE, nDA, DB, SA, SE);
    and (nDA_DB_nSA_SE, nDA, DB, nSA, SE);
    and (nDA_nDB_SA_SE, nDA, nDB, SA, SE);
    and (nDA_nDB_nSA_SE, nDA, nDB, nSA, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SA_int_not, SA_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (DA_check, SA_d, SE_int_not);
  `else
    not  (SA_int_not, SA);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (DA_check, SA, SE_int_not);
  `endif
  buf  (SA_check, SE_int_not);
  and  (DB_check, SA_int_not, SE_int_not);
  or   (CP_check, SI_check, DA_check, SA_check, DB_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    $width (posedge CP &&& DA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFXQD0 (DA, DB, SA, SI, SE, CP, Q);
    input DA, DB, SA, SI, SE, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire DA_d, DB_d, SA_d, SI_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB_d, DA_d, SA_d);
        tsmc_mux (D_i, D, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB, DA, SA);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (DA_DB_SA_SE_SI_SDFCHK, DA_DB_SA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSE_SI_SDFCHK, DA_DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSE_nSI_SDFCHK, DA_DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_SI_SDFCHK, DA_DB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSE_SI_SDFCHK, DA_DB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSE_nSI_SDFCHK, DA_DB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_SI_SDFCHK, DA_nDB_SA_SE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSE_SI_SDFCHK, DA_nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSE_nSI_SDFCHK, DA_nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_SI_SDFCHK, DA_nDB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_SI_SDFCHK, nDA_DB_SA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_SI_SDFCHK, nDA_DB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSE_SI_SDFCHK, nDA_DB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSE_nSI_SDFCHK, nDA_DB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_SI_SDFCHK, nDA_nDB_SA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_SI_SDFCHK, nDA_nDB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_SE_nSI_SDFCHK, DA_DB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_nSI_SDFCHK, DA_DB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_nSI_SDFCHK, DA_nDB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_nSI_SDFCHK, DA_nDB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_nSE_SI_SDFCHK, DA_nDB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_nSE_nSI_SDFCHK, DA_nDB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_nSI_SDFCHK, nDA_DB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_nSE_SI_SDFCHK, nDA_DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_nSE_nSI_SDFCHK, nDA_DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_nSI_SDFCHK, nDA_DB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_nSI_SDFCHK, nDA_nDB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_nSE_SI_SDFCHK, nDA_nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_nSE_nSI_SDFCHK, nDA_nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_nSI_SDFCHK, nDA_nDB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_nSE_SI_SDFCHK, nDA_nDB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_nSE_nSI_SDFCHK, nDA_nDB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DB_SA_nSE_SI_SDFCHK, DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DB_SA_nSE_nSI_SDFCHK, DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDB_SA_nSE_SI_SDFCHK, nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDB_SA_nSE_nSI_SDFCHK, nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nSA_nSE_SI_SDFCHK, DA_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nSA_nSE_nSI_SDFCHK, DA_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nSA_nSE_SI_SDFCHK, nDA_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nSA_nSE_nSI_SDFCHK, nDA_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSE_SI_SDFCHK, DA_nDB_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_nSE_nSI_SDFCHK, DA_nDB_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSE_SI_SDFCHK, nDA_DB_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSE_nSI_SDFCHK, nDA_DB_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SI_SDFCHK, DA_nDB_nSA_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SI_SDFCHK, nDA_DB_SA_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SI_SDFCHK, nDA_nDB_SA_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SI_SDFCHK, nDA_nDB_nSA_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSI_SDFCHK, DA_DB_SA_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSI_SDFCHK, DA_DB_nSA_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSI_SDFCHK, DA_nDB_SA_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSI_SDFCHK, nDA_DB_nSA_nSI, 1'b1);
    tsmc_xbuf (DA_DB_SA_SE_SDFCHK, DA_DB_SA_SE, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_SDFCHK, DA_DB_nSA_SE, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_SDFCHK, DA_nDB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_SDFCHK, nDA_DB_nSA_SE, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_SDFCHK, DA_nDB_nSA_SE, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_SDFCHK, nDA_DB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_SDFCHK, nDA_nDB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_SDFCHK, nDA_nDB_nSA_SE, 1'b1);
  `endif

    not (nDA, DA);
    not (nDB, DB);
    not (nSA, SA);
    not (nSI, SI);
    not (nSE, SE);
    and (DA_DB_SA_SE_SI, DA, DB, SA, SE, SI);
    and (DA_DB_SA_nSE_SI, DA, DB, SA, nSE, SI);
    and (DA_DB_SA_nSE_nSI, DA, DB, SA, nSE, nSI);
    and (DA_DB_nSA_SE_SI, DA, DB, nSA, SE, SI);
    and (DA_DB_nSA_nSE_SI, DA, DB, nSA, nSE, SI);
    and (DA_DB_nSA_nSE_nSI, DA, DB, nSA, nSE, nSI);
    and (DA_nDB_SA_SE_SI, DA, nDB, SA, SE, SI);
    and (DA_nDB_SA_nSE_SI, DA, nDB, SA, nSE, SI);
    and (DA_nDB_SA_nSE_nSI, DA, nDB, SA, nSE, nSI);
    and (DA_nDB_nSA_SE_SI, DA, nDB, nSA, SE, SI);
    and (nDA_DB_SA_SE_SI, nDA, DB, SA, SE, SI);
    and (nDA_DB_nSA_SE_SI, nDA, DB, nSA, SE, SI);
    and (nDA_DB_nSA_nSE_SI, nDA, DB, nSA, nSE, SI);
    and (nDA_DB_nSA_nSE_nSI, nDA, DB, nSA, nSE, nSI);
    and (nDA_nDB_SA_SE_SI, nDA, nDB, SA, SE, SI);
    and (nDA_nDB_nSA_SE_SI, nDA, nDB, nSA, SE, SI);
    and (DA_DB_SA_SE_nSI, DA, DB, SA, SE, nSI);
    and (DA_DB_nSA_SE_nSI, DA, DB, nSA, SE, nSI);
    and (DA_nDB_SA_SE_nSI, DA, nDB, SA, SE, nSI);
    and (DA_nDB_nSA_SE_nSI, DA, nDB, nSA, SE, nSI);
    and (DA_nDB_nSA_nSE_SI, DA, nDB, nSA, nSE, SI);
    and (DA_nDB_nSA_nSE_nSI, DA, nDB, nSA, nSE, nSI);
    and (nDA_DB_SA_SE_nSI, nDA, DB, SA, SE, nSI);
    and (nDA_DB_SA_nSE_SI, nDA, DB, SA, nSE, SI);
    and (nDA_DB_SA_nSE_nSI, nDA, DB, SA, nSE, nSI);
    and (nDA_DB_nSA_SE_nSI, nDA, DB, nSA, SE, nSI);
    and (nDA_nDB_SA_SE_nSI, nDA, nDB, SA, SE, nSI);
    and (nDA_nDB_SA_nSE_SI, nDA, nDB, SA, nSE, SI);
    and (nDA_nDB_SA_nSE_nSI, nDA, nDB, SA, nSE, nSI);
    and (nDA_nDB_nSA_SE_nSI, nDA, nDB, nSA, SE, nSI);
    and (nDA_nDB_nSA_nSE_SI, nDA, nDB, nSA, nSE, SI);
    and (nDA_nDB_nSA_nSE_nSI, nDA, nDB, nSA, nSE, nSI);
    and (DB_SA_nSE_SI, DB, SA, nSE, SI);
    and (DB_SA_nSE_nSI, DB, SA, nSE, nSI);
    and (nDB_SA_nSE_SI, nDB, SA, nSE, SI);
    and (nDB_SA_nSE_nSI, nDB, SA, nSE, nSI);
    and (DA_nSA_nSE_SI, DA, nSA, nSE, SI);
    and (DA_nSA_nSE_nSI, DA, nSA, nSE, nSI);
    and (nDA_nSA_nSE_SI, nDA, nSA, nSE, SI);
    and (nDA_nSA_nSE_nSI, nDA, nSA, nSE, nSI);
    and (DA_nDB_nSE_SI, DA, nDB, nSE, SI);
    and (DA_nDB_nSE_nSI, DA, nDB, nSE, nSI);
    and (nDA_DB_nSE_SI, nDA, DB, nSE, SI);
    and (nDA_DB_nSE_nSI, nDA, DB, nSE, nSI);
    and (DA_nDB_nSA_SI, DA, nDB, nSA, SI);
    and (nDA_DB_SA_SI, nDA, DB, SA, SI);
    and (nDA_nDB_SA_SI, nDA, nDB, SA, SI);
    and (nDA_nDB_nSA_SI, nDA, nDB, nSA, SI);
    and (DA_DB_SA_nSI, DA, DB, SA, nSI);
    and (DA_DB_nSA_nSI, DA, DB, nSA, nSI);
    and (DA_nDB_SA_nSI, DA, nDB, SA, nSI);
    and (nDA_DB_nSA_nSI, nDA, DB, nSA, nSI);
    and (DA_DB_SA_SE, DA, DB, SA, SE);
    and (DA_DB_nSA_SE, DA, DB, nSA, SE);
    and (DA_nDB_SA_SE, DA, nDB, SA, SE);
    and (nDA_DB_nSA_SE, nDA, DB, nSA, SE);
    and (DA_nDB_nSA_SE, DA, nDB, nSA, SE);
    and (nDA_DB_SA_SE, nDA, DB, SA, SE);
    and (nDA_nDB_SA_SE, nDA, nDB, SA, SE);
    and (nDA_nDB_nSA_SE, nDA, nDB, nSA, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SA_int_not, SA_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (DA_check, SA_d, SE_int_not);
  `else
    not  (SA_int_not, SA);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (DA_check, SA, SE_int_not);
  `endif
  buf  (SA_check, SE_int_not);
  and  (DB_check, SA_int_not, SE_int_not);
  or   (CP_check, SI_check, DA_check, SA_check, DB_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    $width (posedge CP &&& DA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFXQD1 (DA, DB, SA, SI, SE, CP, Q);
    input DA, DB, SA, SI, SE, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire DA_d, DB_d, SA_d, SI_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB_d, DA_d, SA_d);
        tsmc_mux (D_i, D, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB, DA, SA);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (DA_DB_SA_SE_SI_SDFCHK, DA_DB_SA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSE_SI_SDFCHK, DA_DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSE_nSI_SDFCHK, DA_DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_SI_SDFCHK, DA_DB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSE_SI_SDFCHK, DA_DB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSE_nSI_SDFCHK, DA_DB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_SI_SDFCHK, DA_nDB_SA_SE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSE_SI_SDFCHK, DA_nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSE_nSI_SDFCHK, DA_nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_SI_SDFCHK, DA_nDB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_SI_SDFCHK, nDA_DB_SA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_SI_SDFCHK, nDA_DB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSE_SI_SDFCHK, nDA_DB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSE_nSI_SDFCHK, nDA_DB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_SI_SDFCHK, nDA_nDB_SA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_SI_SDFCHK, nDA_nDB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_SE_nSI_SDFCHK, DA_DB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_nSI_SDFCHK, DA_DB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_nSI_SDFCHK, DA_nDB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_nSI_SDFCHK, DA_nDB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_nSE_SI_SDFCHK, DA_nDB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_nSE_nSI_SDFCHK, DA_nDB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_nSI_SDFCHK, nDA_DB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_nSE_SI_SDFCHK, nDA_DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_nSE_nSI_SDFCHK, nDA_DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_nSI_SDFCHK, nDA_DB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_nSI_SDFCHK, nDA_nDB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_nSE_SI_SDFCHK, nDA_nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_nSE_nSI_SDFCHK, nDA_nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_nSI_SDFCHK, nDA_nDB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_nSE_SI_SDFCHK, nDA_nDB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_nSE_nSI_SDFCHK, nDA_nDB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DB_SA_nSE_SI_SDFCHK, DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DB_SA_nSE_nSI_SDFCHK, DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDB_SA_nSE_SI_SDFCHK, nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDB_SA_nSE_nSI_SDFCHK, nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nSA_nSE_SI_SDFCHK, DA_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nSA_nSE_nSI_SDFCHK, DA_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nSA_nSE_SI_SDFCHK, nDA_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nSA_nSE_nSI_SDFCHK, nDA_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSE_SI_SDFCHK, DA_nDB_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_nSE_nSI_SDFCHK, DA_nDB_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSE_SI_SDFCHK, nDA_DB_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSE_nSI_SDFCHK, nDA_DB_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SI_SDFCHK, DA_nDB_nSA_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SI_SDFCHK, nDA_DB_SA_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SI_SDFCHK, nDA_nDB_SA_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SI_SDFCHK, nDA_nDB_nSA_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSI_SDFCHK, DA_DB_SA_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSI_SDFCHK, DA_DB_nSA_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSI_SDFCHK, DA_nDB_SA_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSI_SDFCHK, nDA_DB_nSA_nSI, 1'b1);
    tsmc_xbuf (DA_DB_SA_SE_SDFCHK, DA_DB_SA_SE, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_SDFCHK, DA_DB_nSA_SE, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_SDFCHK, DA_nDB_SA_SE, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_SDFCHK, DA_nDB_nSA_SE, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_SDFCHK, nDA_DB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_SDFCHK, nDA_DB_nSA_SE, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_SDFCHK, nDA_nDB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_SDFCHK, nDA_nDB_nSA_SE, 1'b1);
  `endif

    not (nDA, DA);
    not (nDB, DB);
    not (nSA, SA);
    not (nSI, SI);
    not (nSE, SE);
    and (DA_DB_SA_SE_SI, DA, DB, SA, SE, SI);
    and (DA_DB_SA_nSE_SI, DA, DB, SA, nSE, SI);
    and (DA_DB_SA_nSE_nSI, DA, DB, SA, nSE, nSI);
    and (DA_DB_nSA_SE_SI, DA, DB, nSA, SE, SI);
    and (DA_DB_nSA_nSE_SI, DA, DB, nSA, nSE, SI);
    and (DA_DB_nSA_nSE_nSI, DA, DB, nSA, nSE, nSI);
    and (DA_nDB_SA_SE_SI, DA, nDB, SA, SE, SI);
    and (DA_nDB_SA_nSE_SI, DA, nDB, SA, nSE, SI);
    and (DA_nDB_SA_nSE_nSI, DA, nDB, SA, nSE, nSI);
    and (DA_nDB_nSA_SE_SI, DA, nDB, nSA, SE, SI);
    and (nDA_DB_SA_SE_SI, nDA, DB, SA, SE, SI);
    and (nDA_DB_nSA_SE_SI, nDA, DB, nSA, SE, SI);
    and (nDA_DB_nSA_nSE_SI, nDA, DB, nSA, nSE, SI);
    and (nDA_DB_nSA_nSE_nSI, nDA, DB, nSA, nSE, nSI);
    and (nDA_nDB_SA_SE_SI, nDA, nDB, SA, SE, SI);
    and (nDA_nDB_nSA_SE_SI, nDA, nDB, nSA, SE, SI);
    and (DA_DB_SA_SE_nSI, DA, DB, SA, SE, nSI);
    and (DA_DB_nSA_SE_nSI, DA, DB, nSA, SE, nSI);
    and (DA_nDB_SA_SE_nSI, DA, nDB, SA, SE, nSI);
    and (DA_nDB_nSA_SE_nSI, DA, nDB, nSA, SE, nSI);
    and (DA_nDB_nSA_nSE_SI, DA, nDB, nSA, nSE, SI);
    and (DA_nDB_nSA_nSE_nSI, DA, nDB, nSA, nSE, nSI);
    and (nDA_DB_SA_SE_nSI, nDA, DB, SA, SE, nSI);
    and (nDA_DB_SA_nSE_SI, nDA, DB, SA, nSE, SI);
    and (nDA_DB_SA_nSE_nSI, nDA, DB, SA, nSE, nSI);
    and (nDA_DB_nSA_SE_nSI, nDA, DB, nSA, SE, nSI);
    and (nDA_nDB_SA_SE_nSI, nDA, nDB, SA, SE, nSI);
    and (nDA_nDB_SA_nSE_SI, nDA, nDB, SA, nSE, SI);
    and (nDA_nDB_SA_nSE_nSI, nDA, nDB, SA, nSE, nSI);
    and (nDA_nDB_nSA_SE_nSI, nDA, nDB, nSA, SE, nSI);
    and (nDA_nDB_nSA_nSE_SI, nDA, nDB, nSA, nSE, SI);
    and (nDA_nDB_nSA_nSE_nSI, nDA, nDB, nSA, nSE, nSI);
    and (DB_SA_nSE_SI, DB, SA, nSE, SI);
    and (DB_SA_nSE_nSI, DB, SA, nSE, nSI);
    and (nDB_SA_nSE_SI, nDB, SA, nSE, SI);
    and (nDB_SA_nSE_nSI, nDB, SA, nSE, nSI);
    and (DA_nSA_nSE_SI, DA, nSA, nSE, SI);
    and (DA_nSA_nSE_nSI, DA, nSA, nSE, nSI);
    and (nDA_nSA_nSE_SI, nDA, nSA, nSE, SI);
    and (nDA_nSA_nSE_nSI, nDA, nSA, nSE, nSI);
    and (DA_nDB_nSE_SI, DA, nDB, nSE, SI);
    and (DA_nDB_nSE_nSI, DA, nDB, nSE, nSI);
    and (nDA_DB_nSE_SI, nDA, DB, nSE, SI);
    and (nDA_DB_nSE_nSI, nDA, DB, nSE, nSI);
    and (DA_nDB_nSA_SI, DA, nDB, nSA, SI);
    and (nDA_DB_SA_SI, nDA, DB, SA, SI);
    and (nDA_nDB_SA_SI, nDA, nDB, SA, SI);
    and (nDA_nDB_nSA_SI, nDA, nDB, nSA, SI);
    and (DA_DB_SA_nSI, DA, DB, SA, nSI);
    and (DA_DB_nSA_nSI, DA, DB, nSA, nSI);
    and (DA_nDB_SA_nSI, DA, nDB, SA, nSI);
    and (nDA_DB_nSA_nSI, nDA, DB, nSA, nSI);
    and (DA_DB_SA_SE, DA, DB, SA, SE);
    and (DA_DB_nSA_SE, DA, DB, nSA, SE);
    and (DA_nDB_SA_SE, DA, nDB, SA, SE);
    and (DA_nDB_nSA_SE, DA, nDB, nSA, SE);
    and (nDA_DB_SA_SE, nDA, DB, SA, SE);
    and (nDA_DB_nSA_SE, nDA, DB, nSA, SE);
    and (nDA_nDB_SA_SE, nDA, nDB, SA, SE);
    and (nDA_nDB_nSA_SE, nDA, nDB, nSA, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SA_int_not, SA_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (DA_check, SA_d, SE_int_not);
  `else
    not  (SA_int_not, SA);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (DA_check, SA, SE_int_not);
  `endif
  buf  (SA_check, SE_int_not);
  and  (DB_check, SA_int_not, SE_int_not);
  or   (CP_check, SI_check, DA_check, SA_check, DB_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    $width (posedge CP &&& DA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFXQD2 (DA, DB, SA, SI, SE, CP, Q);
    input DA, DB, SA, SI, SE, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire DA_d, DB_d, SA_d, SI_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB_d, DA_d, SA_d);
        tsmc_mux (D_i, D, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB, DA, SA);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (DA_DB_SA_SE_SI_SDFCHK, DA_DB_SA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSE_SI_SDFCHK, DA_DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSE_nSI_SDFCHK, DA_DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_SI_SDFCHK, DA_DB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSE_SI_SDFCHK, DA_DB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSE_nSI_SDFCHK, DA_DB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_SI_SDFCHK, DA_nDB_SA_SE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSE_SI_SDFCHK, DA_nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSE_nSI_SDFCHK, DA_nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_SI_SDFCHK, DA_nDB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_SI_SDFCHK, nDA_DB_SA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_SI_SDFCHK, nDA_DB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSE_SI_SDFCHK, nDA_DB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSE_nSI_SDFCHK, nDA_DB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_SI_SDFCHK, nDA_nDB_SA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_SI_SDFCHK, nDA_nDB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_SE_nSI_SDFCHK, DA_DB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_nSI_SDFCHK, DA_DB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_nSI_SDFCHK, DA_nDB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_nSI_SDFCHK, DA_nDB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_nSE_SI_SDFCHK, DA_nDB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_nSE_nSI_SDFCHK, DA_nDB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_nSI_SDFCHK, nDA_DB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_nSE_SI_SDFCHK, nDA_DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_nSE_nSI_SDFCHK, nDA_DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_nSI_SDFCHK, nDA_DB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_nSI_SDFCHK, nDA_nDB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_nSE_SI_SDFCHK, nDA_nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_nSE_nSI_SDFCHK, nDA_nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_nSI_SDFCHK, nDA_nDB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_nSE_SI_SDFCHK, nDA_nDB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_nSE_nSI_SDFCHK, nDA_nDB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DB_SA_nSE_SI_SDFCHK, DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DB_SA_nSE_nSI_SDFCHK, DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDB_SA_nSE_SI_SDFCHK, nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDB_SA_nSE_nSI_SDFCHK, nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nSA_nSE_SI_SDFCHK, DA_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nSA_nSE_nSI_SDFCHK, DA_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nSA_nSE_SI_SDFCHK, nDA_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nSA_nSE_nSI_SDFCHK, nDA_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSE_SI_SDFCHK, DA_nDB_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_nSE_nSI_SDFCHK, DA_nDB_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSE_SI_SDFCHK, nDA_DB_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSE_nSI_SDFCHK, nDA_DB_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SI_SDFCHK, DA_nDB_nSA_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SI_SDFCHK, nDA_DB_SA_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SI_SDFCHK, nDA_nDB_SA_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SI_SDFCHK, nDA_nDB_nSA_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSI_SDFCHK, DA_DB_SA_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSI_SDFCHK, DA_DB_nSA_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSI_SDFCHK, DA_nDB_SA_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSI_SDFCHK, nDA_DB_nSA_nSI, 1'b1);
    tsmc_xbuf (DA_DB_SA_SE_SDFCHK, DA_DB_SA_SE, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_SDFCHK, DA_DB_nSA_SE, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_SDFCHK, DA_nDB_SA_SE, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_SDFCHK, DA_nDB_nSA_SE, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_SDFCHK, nDA_DB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_SDFCHK, nDA_DB_nSA_SE, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_SDFCHK, nDA_nDB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_SDFCHK, nDA_nDB_nSA_SE, 1'b1);
  `endif

    not (nDA, DA);
    not (nDB, DB);
    not (nSA, SA);
    not (nSI, SI);
    not (nSE, SE);
    and (DA_DB_SA_SE_SI, DA, DB, SA, SE, SI);
    and (DA_DB_SA_nSE_SI, DA, DB, SA, nSE, SI);
    and (DA_DB_SA_nSE_nSI, DA, DB, SA, nSE, nSI);
    and (DA_DB_nSA_SE_SI, DA, DB, nSA, SE, SI);
    and (DA_DB_nSA_nSE_SI, DA, DB, nSA, nSE, SI);
    and (DA_DB_nSA_nSE_nSI, DA, DB, nSA, nSE, nSI);
    and (DA_nDB_SA_SE_SI, DA, nDB, SA, SE, SI);
    and (DA_nDB_SA_nSE_SI, DA, nDB, SA, nSE, SI);
    and (DA_nDB_SA_nSE_nSI, DA, nDB, SA, nSE, nSI);
    and (DA_nDB_nSA_SE_SI, DA, nDB, nSA, SE, SI);
    and (nDA_DB_SA_SE_SI, nDA, DB, SA, SE, SI);
    and (nDA_DB_nSA_SE_SI, nDA, DB, nSA, SE, SI);
    and (nDA_DB_nSA_nSE_SI, nDA, DB, nSA, nSE, SI);
    and (nDA_DB_nSA_nSE_nSI, nDA, DB, nSA, nSE, nSI);
    and (nDA_nDB_SA_SE_SI, nDA, nDB, SA, SE, SI);
    and (nDA_nDB_nSA_SE_SI, nDA, nDB, nSA, SE, SI);
    and (DA_DB_SA_SE_nSI, DA, DB, SA, SE, nSI);
    and (DA_DB_nSA_SE_nSI, DA, DB, nSA, SE, nSI);
    and (DA_nDB_SA_SE_nSI, DA, nDB, SA, SE, nSI);
    and (DA_nDB_nSA_SE_nSI, DA, nDB, nSA, SE, nSI);
    and (DA_nDB_nSA_nSE_SI, DA, nDB, nSA, nSE, SI);
    and (DA_nDB_nSA_nSE_nSI, DA, nDB, nSA, nSE, nSI);
    and (nDA_DB_SA_SE_nSI, nDA, DB, SA, SE, nSI);
    and (nDA_DB_SA_nSE_SI, nDA, DB, SA, nSE, SI);
    and (nDA_DB_SA_nSE_nSI, nDA, DB, SA, nSE, nSI);
    and (nDA_DB_nSA_SE_nSI, nDA, DB, nSA, SE, nSI);
    and (nDA_nDB_SA_SE_nSI, nDA, nDB, SA, SE, nSI);
    and (nDA_nDB_SA_nSE_SI, nDA, nDB, SA, nSE, SI);
    and (nDA_nDB_SA_nSE_nSI, nDA, nDB, SA, nSE, nSI);
    and (nDA_nDB_nSA_SE_nSI, nDA, nDB, nSA, SE, nSI);
    and (nDA_nDB_nSA_nSE_SI, nDA, nDB, nSA, nSE, SI);
    and (nDA_nDB_nSA_nSE_nSI, nDA, nDB, nSA, nSE, nSI);
    and (DB_SA_nSE_SI, DB, SA, nSE, SI);
    and (DB_SA_nSE_nSI, DB, SA, nSE, nSI);
    and (nDB_SA_nSE_SI, nDB, SA, nSE, SI);
    and (nDB_SA_nSE_nSI, nDB, SA, nSE, nSI);
    and (DA_nSA_nSE_SI, DA, nSA, nSE, SI);
    and (DA_nSA_nSE_nSI, DA, nSA, nSE, nSI);
    and (nDA_nSA_nSE_SI, nDA, nSA, nSE, SI);
    and (nDA_nSA_nSE_nSI, nDA, nSA, nSE, nSI);
    and (DA_nDB_nSE_SI, DA, nDB, nSE, SI);
    and (DA_nDB_nSE_nSI, DA, nDB, nSE, nSI);
    and (nDA_DB_nSE_SI, nDA, DB, nSE, SI);
    and (nDA_DB_nSE_nSI, nDA, DB, nSE, nSI);
    and (DA_nDB_nSA_SI, DA, nDB, nSA, SI);
    and (nDA_DB_SA_SI, nDA, DB, SA, SI);
    and (nDA_nDB_SA_SI, nDA, nDB, SA, SI);
    and (nDA_nDB_nSA_SI, nDA, nDB, nSA, SI);
    and (DA_DB_SA_nSI, DA, DB, SA, nSI);
    and (DA_DB_nSA_nSI, DA, DB, nSA, nSI);
    and (DA_nDB_SA_nSI, DA, nDB, SA, nSI);
    and (nDA_DB_nSA_nSI, nDA, DB, nSA, nSI);
    and (DA_DB_SA_SE, DA, DB, SA, SE);
    and (DA_DB_nSA_SE, DA, DB, nSA, SE);
    and (DA_nDB_SA_SE, DA, nDB, SA, SE);
    and (DA_nDB_nSA_SE, DA, nDB, nSA, SE);
    and (nDA_DB_SA_SE, nDA, DB, SA, SE);
    and (nDA_DB_nSA_SE, nDA, DB, nSA, SE);
    and (nDA_nDB_SA_SE, nDA, nDB, SA, SE);
    and (nDA_nDB_nSA_SE, nDA, nDB, nSA, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SA_int_not, SA_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (DA_check, SA_d, SE_int_not);
  `else
    not  (SA_int_not, SA);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (DA_check, SA, SE_int_not);
  `endif
  buf  (SA_check, SE_int_not);
  and  (DB_check, SA_int_not, SE_int_not);
  or   (CP_check, SI_check, DA_check, SA_check, DB_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    $width (posedge CP &&& DA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFXQD4 (DA, DB, SA, SI, SE, CP, Q);
    input DA, DB, SA, SI, SE, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire DA_d, DB_d, SA_d, SI_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB_d, DA_d, SA_d);
        tsmc_mux (D_i, D, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB, DA, SA);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (DA_DB_SA_SE_SI_SDFCHK, DA_DB_SA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSE_SI_SDFCHK, DA_DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSE_nSI_SDFCHK, DA_DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_SI_SDFCHK, DA_DB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSE_SI_SDFCHK, DA_DB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSE_nSI_SDFCHK, DA_DB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_SI_SDFCHK, DA_nDB_SA_SE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSE_SI_SDFCHK, DA_nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSE_nSI_SDFCHK, DA_nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_SI_SDFCHK, DA_nDB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_SI_SDFCHK, nDA_DB_SA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_SI_SDFCHK, nDA_DB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSE_SI_SDFCHK, nDA_DB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSE_nSI_SDFCHK, nDA_DB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_SI_SDFCHK, nDA_nDB_SA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_SI_SDFCHK, nDA_nDB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_SE_nSI_SDFCHK, DA_DB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_nSI_SDFCHK, DA_DB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_nSI_SDFCHK, DA_nDB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_nSI_SDFCHK, DA_nDB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_nSE_SI_SDFCHK, DA_nDB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_nSE_nSI_SDFCHK, DA_nDB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_nSI_SDFCHK, nDA_DB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_nSE_SI_SDFCHK, nDA_DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_nSE_nSI_SDFCHK, nDA_DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_nSI_SDFCHK, nDA_DB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_nSI_SDFCHK, nDA_nDB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_nSE_SI_SDFCHK, nDA_nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_nSE_nSI_SDFCHK, nDA_nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_nSI_SDFCHK, nDA_nDB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_nSE_SI_SDFCHK, nDA_nDB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_nSE_nSI_SDFCHK, nDA_nDB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DB_SA_nSE_SI_SDFCHK, DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DB_SA_nSE_nSI_SDFCHK, DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDB_SA_nSE_SI_SDFCHK, nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDB_SA_nSE_nSI_SDFCHK, nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nSA_nSE_SI_SDFCHK, DA_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nSA_nSE_nSI_SDFCHK, DA_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nSA_nSE_SI_SDFCHK, nDA_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nSA_nSE_nSI_SDFCHK, nDA_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSE_SI_SDFCHK, DA_nDB_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_nSE_nSI_SDFCHK, DA_nDB_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSE_SI_SDFCHK, nDA_DB_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSE_nSI_SDFCHK, nDA_DB_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SI_SDFCHK, DA_nDB_nSA_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SI_SDFCHK, nDA_DB_SA_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SI_SDFCHK, nDA_nDB_SA_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SI_SDFCHK, nDA_nDB_nSA_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSI_SDFCHK, DA_DB_SA_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSI_SDFCHK, DA_DB_nSA_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSI_SDFCHK, DA_nDB_SA_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSI_SDFCHK, nDA_DB_nSA_nSI, 1'b1);
    tsmc_xbuf (DA_DB_SA_SE_SDFCHK, DA_DB_SA_SE, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_SDFCHK, DA_DB_nSA_SE, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_SDFCHK, DA_nDB_SA_SE, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_SDFCHK, DA_nDB_nSA_SE, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_SDFCHK, nDA_DB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_SDFCHK, nDA_DB_nSA_SE, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_SDFCHK, nDA_nDB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_SDFCHK, nDA_nDB_nSA_SE, 1'b1);
  `endif

    not (nDA, DA);
    not (nDB, DB);
    not (nSA, SA);
    not (nSI, SI);
    not (nSE, SE);
    and (DA_DB_SA_SE_SI, DA, DB, SA, SE, SI);
    and (DA_DB_SA_nSE_SI, DA, DB, SA, nSE, SI);
    and (DA_DB_SA_nSE_nSI, DA, DB, SA, nSE, nSI);
    and (DA_DB_nSA_SE_SI, DA, DB, nSA, SE, SI);
    and (DA_DB_nSA_nSE_SI, DA, DB, nSA, nSE, SI);
    and (DA_DB_nSA_nSE_nSI, DA, DB, nSA, nSE, nSI);
    and (DA_nDB_SA_SE_SI, DA, nDB, SA, SE, SI);
    and (DA_nDB_SA_nSE_SI, DA, nDB, SA, nSE, SI);
    and (DA_nDB_SA_nSE_nSI, DA, nDB, SA, nSE, nSI);
    and (DA_nDB_nSA_SE_SI, DA, nDB, nSA, SE, SI);
    and (nDA_DB_SA_SE_SI, nDA, DB, SA, SE, SI);
    and (nDA_DB_nSA_SE_SI, nDA, DB, nSA, SE, SI);
    and (nDA_DB_nSA_nSE_SI, nDA, DB, nSA, nSE, SI);
    and (nDA_DB_nSA_nSE_nSI, nDA, DB, nSA, nSE, nSI);
    and (nDA_nDB_SA_SE_SI, nDA, nDB, SA, SE, SI);
    and (nDA_nDB_nSA_SE_SI, nDA, nDB, nSA, SE, SI);
    and (DA_DB_SA_SE_nSI, DA, DB, SA, SE, nSI);
    and (DA_DB_nSA_SE_nSI, DA, DB, nSA, SE, nSI);
    and (DA_nDB_SA_SE_nSI, DA, nDB, SA, SE, nSI);
    and (DA_nDB_nSA_SE_nSI, DA, nDB, nSA, SE, nSI);
    and (DA_nDB_nSA_nSE_SI, DA, nDB, nSA, nSE, SI);
    and (DA_nDB_nSA_nSE_nSI, DA, nDB, nSA, nSE, nSI);
    and (nDA_DB_SA_SE_nSI, nDA, DB, SA, SE, nSI);
    and (nDA_DB_SA_nSE_SI, nDA, DB, SA, nSE, SI);
    and (nDA_DB_SA_nSE_nSI, nDA, DB, SA, nSE, nSI);
    and (nDA_DB_nSA_SE_nSI, nDA, DB, nSA, SE, nSI);
    and (nDA_nDB_SA_SE_nSI, nDA, nDB, SA, SE, nSI);
    and (nDA_nDB_SA_nSE_SI, nDA, nDB, SA, nSE, SI);
    and (nDA_nDB_SA_nSE_nSI, nDA, nDB, SA, nSE, nSI);
    and (nDA_nDB_nSA_SE_nSI, nDA, nDB, nSA, SE, nSI);
    and (nDA_nDB_nSA_nSE_SI, nDA, nDB, nSA, nSE, SI);
    and (nDA_nDB_nSA_nSE_nSI, nDA, nDB, nSA, nSE, nSI);
    and (DB_SA_nSE_SI, DB, SA, nSE, SI);
    and (DB_SA_nSE_nSI, DB, SA, nSE, nSI);
    and (nDB_SA_nSE_SI, nDB, SA, nSE, SI);
    and (nDB_SA_nSE_nSI, nDB, SA, nSE, nSI);
    and (DA_nSA_nSE_SI, DA, nSA, nSE, SI);
    and (DA_nSA_nSE_nSI, DA, nSA, nSE, nSI);
    and (nDA_nSA_nSE_SI, nDA, nSA, nSE, SI);
    and (nDA_nSA_nSE_nSI, nDA, nSA, nSE, nSI);
    and (DA_nDB_nSE_SI, DA, nDB, nSE, SI);
    and (DA_nDB_nSE_nSI, DA, nDB, nSE, nSI);
    and (nDA_DB_nSE_SI, nDA, DB, nSE, SI);
    and (nDA_DB_nSE_nSI, nDA, DB, nSE, nSI);
    and (DA_nDB_nSA_SI, DA, nDB, nSA, SI);
    and (nDA_DB_SA_SI, nDA, DB, SA, SI);
    and (nDA_nDB_SA_SI, nDA, nDB, SA, SI);
    and (nDA_nDB_nSA_SI, nDA, nDB, nSA, SI);
    and (DA_DB_SA_nSI, DA, DB, SA, nSI);
    and (DA_DB_nSA_nSI, DA, DB, nSA, nSI);
    and (DA_nDB_SA_nSI, DA, nDB, SA, nSI);
    and (nDA_DB_nSA_nSI, nDA, DB, nSA, nSI);
    and (DA_DB_SA_SE, DA, DB, SA, SE);
    and (DA_DB_nSA_SE, DA, DB, nSA, SE);
    and (DA_nDB_SA_SE, DA, nDB, SA, SE);
    and (DA_nDB_nSA_SE, DA, nDB, nSA, SE);
    and (nDA_DB_SA_SE, nDA, DB, SA, SE);
    and (nDA_DB_nSA_SE, nDA, DB, nSA, SE);
    and (nDA_nDB_SA_SE, nDA, nDB, SA, SE);
    and (nDA_nDB_nSA_SE, nDA, nDB, nSA, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SA_int_not, SA_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (DA_check, SA_d, SE_int_not);
  `else
    not  (SA_int_not, SA);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (DA_check, SA, SE_int_not);
  `endif
  buf  (SA_check, SE_int_not);
  and  (DB_check, SA_int_not, SE_int_not);
  or   (CP_check, SI_check, DA_check, SA_check, DB_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    $width (posedge CP &&& DA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDF4CQD0 (E, SE, CP, SI, D, Q);
    input E, SE, CP, SI, D;
    output Q;
    reg notifier;
    `ifdef NTC
        wire E_d, SE_d, CP_d, SI_d, D_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_E_SE_SI_SDFCHK, D_E_SE_SI, 1'b1);
    tsmc_xbuf (D_nE_SE_SI_SDFCHK, D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nD_E_SE_SI_SDFCHK, nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SE_SI_SDFCHK, nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_SI_SDFCHK, D_E_nSE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_nSI_SDFCHK, D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_E_SE_nSI_SDFCHK, D_E_SE_nSI, 1'b1);
    tsmc_xbuf (D_nE_SE_nSI_SDFCHK, D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nD_E_SE_nSI_SDFCHK, nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_SE_nSI_SDFCHK, nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nD_E_nSE_SI_SDFCHK, nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (nD_E_nSE_nSI_SDFCHK, nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (E_nSE_SI_SDFCHK, E_nSE_SI, 1'b1);
    tsmc_xbuf (E_nSE_nSI_SDFCHK, E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nE_SI_SDFCHK, D_nE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SI_SDFCHK, nD_nE_SI, 1'b1);
    tsmc_xbuf (nD_E_SI_SDFCHK, nD_E_SI, 1'b1);
    tsmc_xbuf (D_E_nSI_SDFCHK, D_E_nSI, 1'b1);
    tsmc_xbuf (D_nE_nSI_SDFCHK, D_nE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_nSI_SDFCHK, nD_nE_nSI, 1'b1);
    tsmc_xbuf (D_E_SE_SDFCHK, D_E_SE, 1'b1);
    tsmc_xbuf (nD_E_SE_SDFCHK, nD_E_SE, 1'b1);
    tsmc_xbuf (D_nE_SE_SDFCHK, D_nE_SE, 1'b1);
    tsmc_xbuf (nD_nE_SE_SDFCHK, nD_nE_SE, 1'b1);
  `endif

    not (nE, E);
    not (nSE, SE);
    not (nSI, SI);
    not (nD, D);
    and (D_E_SE_SI, D, E, SE, SI);
    and (D_nE_SE_SI, D, nE, SE, SI);
    and (nD_E_SE_SI, nD, E, SE, SI);
    and (nD_nE_SE_SI, nD, nE, SE, SI);
    and (D_E_nSE_SI, D, E, nSE, SI);
    and (D_E_nSE_nSI, D, E, nSE, nSI);
    and (D_E_SE_nSI, D, E, SE, nSI);
    and (D_nE_SE_nSI, D, nE, SE, nSI);
    and (nD_E_SE_nSI, nD, E, SE, nSI);
    and (nD_nE_SE_nSI, nD, nE, SE, nSI);
    and (nD_E_nSE_SI, nD, E, nSE, SI);
    and (nD_E_nSE_nSI, nD, E, nSE, nSI);
    and (E_nSE_SI, E, nSE, SI);
    and (E_nSE_nSI, E, nSE, nSI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (D_nE_SI, D, nE, SI);
    and (nD_nE_SI, nD, nE, SI);
    and (nD_E_SI, nD, E, SI);
    and (D_E_nSI, D, E, nSI);
    and (D_nE_nSI, D, nE, nSI);
    and (nD_nE_nSI, nD, nE, nSI);
    and (D_E_SE, D, E, SE);
    and (nD_E_SE, nD, E, SE);
    and (D_nE_SE, D, nE, SE);
    and (nD_nE_SE, nD, nE, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDF4CQD1 (E, SE, CP, SI, D, Q);
    input E, SE, CP, SI, D;
    output Q;
    reg notifier;
    `ifdef NTC
        wire E_d, SE_d, CP_d, SI_d, D_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_E_SE_SI_SDFCHK, D_E_SE_SI, 1'b1);
    tsmc_xbuf (D_nE_SE_SI_SDFCHK, D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nD_E_SE_SI_SDFCHK, nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SE_SI_SDFCHK, nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_SI_SDFCHK, D_E_nSE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_nSI_SDFCHK, D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_E_SE_nSI_SDFCHK, D_E_SE_nSI, 1'b1);
    tsmc_xbuf (D_nE_SE_nSI_SDFCHK, D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nD_E_SE_nSI_SDFCHK, nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_SE_nSI_SDFCHK, nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nD_E_nSE_SI_SDFCHK, nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (nD_E_nSE_nSI_SDFCHK, nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (E_nSE_SI_SDFCHK, E_nSE_SI, 1'b1);
    tsmc_xbuf (E_nSE_nSI_SDFCHK, E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nE_SI_SDFCHK, D_nE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SI_SDFCHK, nD_nE_SI, 1'b1);
    tsmc_xbuf (nD_E_SI_SDFCHK, nD_E_SI, 1'b1);
    tsmc_xbuf (D_E_nSI_SDFCHK, D_E_nSI, 1'b1);
    tsmc_xbuf (D_nE_nSI_SDFCHK, D_nE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_nSI_SDFCHK, nD_nE_nSI, 1'b1);
    tsmc_xbuf (D_E_SE_SDFCHK, D_E_SE, 1'b1);
    tsmc_xbuf (nD_E_SE_SDFCHK, nD_E_SE, 1'b1);
    tsmc_xbuf (D_nE_SE_SDFCHK, D_nE_SE, 1'b1);
    tsmc_xbuf (nD_nE_SE_SDFCHK, nD_nE_SE, 1'b1);
  `endif

    not (nE, E);
    not (nSE, SE);
    not (nSI, SI);
    not (nD, D);
    and (D_E_SE_SI, D, E, SE, SI);
    and (D_nE_SE_SI, D, nE, SE, SI);
    and (nD_E_SE_SI, nD, E, SE, SI);
    and (nD_nE_SE_SI, nD, nE, SE, SI);
    and (D_E_nSE_SI, D, E, nSE, SI);
    and (D_E_nSE_nSI, D, E, nSE, nSI);
    and (D_E_SE_nSI, D, E, SE, nSI);
    and (D_nE_SE_nSI, D, nE, SE, nSI);
    and (nD_E_SE_nSI, nD, E, SE, nSI);
    and (nD_nE_SE_nSI, nD, nE, SE, nSI);
    and (nD_E_nSE_SI, nD, E, nSE, SI);
    and (nD_E_nSE_nSI, nD, E, nSE, nSI);
    and (E_nSE_SI, E, nSE, SI);
    and (E_nSE_nSI, E, nSE, nSI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (D_nE_SI, D, nE, SI);
    and (nD_nE_SI, nD, nE, SI);
    and (nD_E_SI, nD, E, SI);
    and (D_E_nSI, D, E, nSI);
    and (D_nE_nSI, D, nE, nSI);
    and (nD_nE_nSI, nD, nE, nSI);
    and (D_E_SE, D, E, SE);
    and (nD_E_SE, nD, E, SE);
    and (D_nE_SE, D, nE, SE);
    and (nD_nE_SE, nD, nE, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDF4CQD2 (E, SE, CP, SI, D, Q);
    input E, SE, CP, SI, D;
    output Q;
    reg notifier;
    `ifdef NTC
        wire E_d, SE_d, CP_d, SI_d, D_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_E_SE_SI_SDFCHK, D_E_SE_SI, 1'b1);
    tsmc_xbuf (D_nE_SE_SI_SDFCHK, D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nD_E_SE_SI_SDFCHK, nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SE_SI_SDFCHK, nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_SI_SDFCHK, D_E_nSE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_nSI_SDFCHK, D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_E_SE_nSI_SDFCHK, D_E_SE_nSI, 1'b1);
    tsmc_xbuf (D_nE_SE_nSI_SDFCHK, D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nD_E_SE_nSI_SDFCHK, nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_SE_nSI_SDFCHK, nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nD_E_nSE_SI_SDFCHK, nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (nD_E_nSE_nSI_SDFCHK, nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (E_nSE_SI_SDFCHK, E_nSE_SI, 1'b1);
    tsmc_xbuf (E_nSE_nSI_SDFCHK, E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nE_SI_SDFCHK, D_nE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SI_SDFCHK, nD_nE_SI, 1'b1);
    tsmc_xbuf (nD_E_SI_SDFCHK, nD_E_SI, 1'b1);
    tsmc_xbuf (D_E_nSI_SDFCHK, D_E_nSI, 1'b1);
    tsmc_xbuf (D_nE_nSI_SDFCHK, D_nE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_nSI_SDFCHK, nD_nE_nSI, 1'b1);
    tsmc_xbuf (D_E_SE_SDFCHK, D_E_SE, 1'b1);
    tsmc_xbuf (nD_E_SE_SDFCHK, nD_E_SE, 1'b1);
    tsmc_xbuf (D_nE_SE_SDFCHK, D_nE_SE, 1'b1);
    tsmc_xbuf (nD_nE_SE_SDFCHK, nD_nE_SE, 1'b1);
  `endif

    not (nE, E);
    not (nSE, SE);
    not (nSI, SI);
    not (nD, D);
    and (D_E_SE_SI, D, E, SE, SI);
    and (D_nE_SE_SI, D, nE, SE, SI);
    and (nD_E_SE_SI, nD, E, SE, SI);
    and (nD_nE_SE_SI, nD, nE, SE, SI);
    and (D_E_nSE_SI, D, E, nSE, SI);
    and (D_E_nSE_nSI, D, E, nSE, nSI);
    and (D_E_SE_nSI, D, E, SE, nSI);
    and (D_nE_SE_nSI, D, nE, SE, nSI);
    and (nD_E_SE_nSI, nD, E, SE, nSI);
    and (nD_nE_SE_nSI, nD, nE, SE, nSI);
    and (nD_E_nSE_SI, nD, E, nSE, SI);
    and (nD_E_nSE_nSI, nD, E, nSE, nSI);
    and (E_nSE_SI, E, nSE, SI);
    and (E_nSE_nSI, E, nSE, nSI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (D_nE_SI, D, nE, SI);
    and (nD_nE_SI, nD, nE, SI);
    and (nD_E_SI, nD, E, SI);
    and (D_E_nSI, D, E, nSI);
    and (D_nE_nSI, D, nE, nSI);
    and (nD_nE_nSI, nD, nE, nSI);
    and (D_E_SE, D, E, SE);
    and (nD_E_SE, nD, E, SE);
    and (D_nE_SE, D, nE, SE);
    and (nD_nE_SE, nD, nE, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDF4CQD4 (E, SE, CP, SI, D, Q);
    input E, SE, CP, SI, D;
    output Q;
    reg notifier;
    `ifdef NTC
        wire E_d, SE_d, CP_d, SI_d, D_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_E_SE_SI_SDFCHK, D_E_SE_SI, 1'b1);
    tsmc_xbuf (D_nE_SE_SI_SDFCHK, D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nD_E_SE_SI_SDFCHK, nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SE_SI_SDFCHK, nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_SI_SDFCHK, D_E_nSE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_nSI_SDFCHK, D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_E_SE_nSI_SDFCHK, D_E_SE_nSI, 1'b1);
    tsmc_xbuf (D_nE_SE_nSI_SDFCHK, D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nD_E_SE_nSI_SDFCHK, nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_SE_nSI_SDFCHK, nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nD_E_nSE_SI_SDFCHK, nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (nD_E_nSE_nSI_SDFCHK, nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (E_nSE_SI_SDFCHK, E_nSE_SI, 1'b1);
    tsmc_xbuf (E_nSE_nSI_SDFCHK, E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nE_SI_SDFCHK, D_nE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SI_SDFCHK, nD_nE_SI, 1'b1);
    tsmc_xbuf (nD_E_SI_SDFCHK, nD_E_SI, 1'b1);
    tsmc_xbuf (D_E_nSI_SDFCHK, D_E_nSI, 1'b1);
    tsmc_xbuf (D_nE_nSI_SDFCHK, D_nE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_nSI_SDFCHK, nD_nE_nSI, 1'b1);
    tsmc_xbuf (D_E_SE_SDFCHK, D_E_SE, 1'b1);
    tsmc_xbuf (nD_E_SE_SDFCHK, nD_E_SE, 1'b1);
    tsmc_xbuf (D_nE_SE_SDFCHK, D_nE_SE, 1'b1);
    tsmc_xbuf (nD_nE_SE_SDFCHK, nD_nE_SE, 1'b1);
  `endif

    not (nE, E);
    not (nSE, SE);
    not (nSI, SI);
    not (nD, D);
    and (D_E_SE_SI, D, E, SE, SI);
    and (D_nE_SE_SI, D, nE, SE, SI);
    and (nD_E_SE_SI, nD, E, SE, SI);
    and (nD_nE_SE_SI, nD, nE, SE, SI);
    and (D_E_nSE_SI, D, E, nSE, SI);
    and (D_E_nSE_nSI, D, E, nSE, nSI);
    and (D_E_SE_nSI, D, E, SE, nSI);
    and (D_nE_SE_nSI, D, nE, SE, nSI);
    and (nD_E_SE_nSI, nD, E, SE, nSI);
    and (nD_nE_SE_nSI, nD, nE, SE, nSI);
    and (nD_E_nSE_SI, nD, E, nSE, SI);
    and (nD_E_nSE_nSI, nD, E, nSE, nSI);
    and (E_nSE_SI, E, nSE, SI);
    and (E_nSE_nSI, E, nSE, nSI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (D_nE_SI, D, nE, SI);
    and (nD_nE_SI, nD, nE, SI);
    and (nD_E_SI, nD, E, SI);
    and (D_E_nSI, D, E, nSI);
    and (D_nE_nSI, D, nE, nSI);
    and (nD_nE_nSI, nD, nE, nSI);
    and (D_E_SE, D, E, SE);
    and (nD_E_SE, nD, E, SE);
    and (D_nE_SE, D, nE, SE);
    and (nD_nE_SE, nD, nE, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFCND0 (E, SE, CP, SI, D, CDN, Q, QN);
    input E, SE, CP, SI, D, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire E_d, SE_d, CP_d, SI_d, D_d;
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_E_SE_SI_SDFCHK, CP_D_E_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_E_SE_nSI_SDFCHK, CP_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_E_nSE_SI_SDFCHK, CP_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_E_nSE_nSI_SDFCHK, CP_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_E_SE_SI_SDFCHK, CP_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_E_SE_nSI_SDFCHK, CP_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_E_nSE_SI_SDFCHK, CP_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_E_nSE_nSI_SDFCHK, CP_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nE_SE_SI_SDFCHK, CP_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_nE_SE_nSI_SDFCHK, CP_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nE_nSE_SI_SDFCHK, CP_D_nE_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nE_nSE_nSI_SDFCHK, CP_D_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nE_SE_SI_SDFCHK, CP_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nE_SE_nSI_SDFCHK, CP_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nE_nSE_SI_SDFCHK, CP_nD_nE_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nE_nSE_nSI_SDFCHK, CP_nD_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_E_SE_SI_SDFCHK, nCP_D_E_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_E_SE_nSI_SDFCHK, nCP_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_E_nSE_SI_SDFCHK, nCP_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_E_nSE_nSI_SDFCHK, nCP_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_E_SE_SI_SDFCHK, nCP_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_E_SE_nSI_SDFCHK, nCP_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_E_nSE_SI_SDFCHK, nCP_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_E_nSE_nSI_SDFCHK, nCP_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nE_SE_SI_SDFCHK, nCP_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nE_SE_nSI_SDFCHK, nCP_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nE_nSE_SI_SDFCHK, nCP_D_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nE_nSE_nSI_SDFCHK, nCP_D_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nE_SE_SI_SDFCHK, nCP_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nE_SE_nSI_SDFCHK, nCP_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nE_nSE_SI_SDFCHK, nCP_nD_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nE_nSE_nSI_SDFCHK, nCP_nD_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_E_SE_SI_SDFCHK, CDN_D_E_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_E_nSE_SI_SDFCHK, CDN_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_E_nSE_nSI_SDFCHK, CDN_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_E_SE_SI_SDFCHK, CDN_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nE_SE_SI_SDFCHK, CDN_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SE_SI_SDFCHK, CDN_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_E_SE_nSI_SDFCHK, CDN_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_E_SE_nSI_SDFCHK, CDN_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_E_nSE_SI_SDFCHK, CDN_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_E_nSE_nSI_SDFCHK, CDN_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_nE_SE_nSI_SDFCHK, CDN_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SE_nSI_SDFCHK, CDN_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_E_nSE_SI_SDFCHK, CDN_E_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_E_nSE_nSI_SDFCHK, CDN_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_nE_SI_SDFCHK, CDN_D_nE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SI_SDFCHK, CDN_nD_nE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_E_SI_SDFCHK, CDN_nD_E_SI, 1'b1);
    tsmc_xbuf (CDN_D_E_nSI_SDFCHK, CDN_D_E_nSI, 1'b1);
    tsmc_xbuf (CDN_D_nE_nSI_SDFCHK, CDN_D_nE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nE_nSI_SDFCHK, CDN_nD_nE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_E_SE_SDFCHK, CDN_D_E_SE, 1'b1);
    tsmc_xbuf (CDN_D_nE_SE_SDFCHK, CDN_D_nE_SE, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SE_SDFCHK, CDN_nD_nE_SE, 1'b1);
    tsmc_xbuf (CDN_nD_E_SE_SDFCHK, CDN_nD_E_SE, 1'b1);
    tsmc_xbuf (D_E_SE_SI_SDFCHK, D_E_SE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_SI_SDFCHK, D_E_nSE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_nSI_SDFCHK, D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_E_SE_SI_SDFCHK, nD_E_SE_SI, 1'b1);
    tsmc_xbuf (D_nE_SE_SI_SDFCHK, D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SE_SI_SDFCHK, nD_nE_SE_SI, 1'b1);
  `endif

    not (nE, E);
    not (nSE, SE);
    not (nCP, CP);
    not (nSI, SI);
    not (nD, D);
    and (CP_D_E_SE_SI, CP, D, E, SE, SI);
    and (CP_D_E_SE_nSI, CP, D, E, SE, nSI);
    and (CP_D_E_nSE_SI, CP, D, E, nSE, SI);
    and (CP_D_E_nSE_nSI, CP, D, E, nSE, nSI);
    and (CP_nD_E_SE_SI, CP, nD, E, SE, SI);
    and (CP_nD_E_SE_nSI, CP, nD, E, SE, nSI);
    and (CP_nD_E_nSE_SI, CP, nD, E, nSE, SI);
    and (CP_nD_E_nSE_nSI, CP, nD, E, nSE, nSI);
    and (CP_D_nE_SE_SI, CP, D, nE, SE, SI);
    and (CP_D_nE_SE_nSI, CP, D, nE, SE, nSI);
    and (CP_D_nE_nSE_SI, CP, D, nE, nSE, SI);
    and (CP_D_nE_nSE_nSI, CP, D, nE, nSE, nSI);
    and (CP_nD_nE_SE_SI, CP, nD, nE, SE, SI);
    and (CP_nD_nE_SE_nSI, CP, nD, nE, SE, nSI);
    and (CP_nD_nE_nSE_SI, CP, nD, nE, nSE, SI);
    and (CP_nD_nE_nSE_nSI, CP, nD, nE, nSE, nSI);
    and (nCP_D_E_SE_SI, nCP, D, E, SE, SI);
    and (nCP_D_E_SE_nSI, nCP, D, E, SE, nSI);
    and (nCP_D_E_nSE_SI, nCP, D, E, nSE, SI);
    and (nCP_D_E_nSE_nSI, nCP, D, E, nSE, nSI);
    and (nCP_nD_E_SE_SI, nCP, nD, E, SE, SI);
    and (nCP_nD_E_SE_nSI, nCP, nD, E, SE, nSI);
    and (nCP_nD_E_nSE_SI, nCP, nD, E, nSE, SI);
    and (nCP_nD_E_nSE_nSI, nCP, nD, E, nSE, nSI);
    and (nCP_D_nE_SE_SI, nCP, D, nE, SE, SI);
    and (nCP_D_nE_SE_nSI, nCP, D, nE, SE, nSI);
    and (nCP_D_nE_nSE_SI, nCP, D, nE, nSE, SI);
    and (nCP_D_nE_nSE_nSI, nCP, D, nE, nSE, nSI);
    and (nCP_nD_nE_SE_SI, nCP, nD, nE, SE, SI);
    and (nCP_nD_nE_SE_nSI, nCP, nD, nE, SE, nSI);
    and (nCP_nD_nE_nSE_SI, nCP, nD, nE, nSE, SI);
    and (nCP_nD_nE_nSE_nSI, nCP, nD, nE, nSE, nSI);
    and (CDN_D_E_SE_SI, CDN, D, E, SE, SI);
    and (CDN_D_E_nSE_SI, CDN, D, E, nSE, SI);
    and (CDN_D_E_nSE_nSI, CDN, D, E, nSE, nSI);
    and (CDN_nD_E_SE_SI, CDN, nD, E, SE, SI);
    and (CDN_D_nE_SE_SI, CDN, D, nE, SE, SI);
    and (CDN_nD_nE_SE_SI, CDN, nD, nE, SE, SI);
    and (CDN_D_E_SE_nSI, CDN, D, E, SE, nSI);
    and (CDN_nD_E_SE_nSI, CDN, nD, E, SE, nSI);
    and (CDN_nD_E_nSE_SI, CDN, nD, E, nSE, SI);
    and (CDN_nD_E_nSE_nSI, CDN, nD, E, nSE, nSI);
    and (CDN_D_nE_SE_nSI, CDN, D, nE, SE, nSI);
    and (CDN_nD_nE_SE_nSI, CDN, nD, nE, SE, nSI);
    and (CDN_E_nSE_SI, CDN, E, nSE, SI);
    and (CDN_E_nSE_nSI, CDN, E, nSE, nSI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_D_nE_SI, CDN, D, nE, SI);
    and (CDN_nD_nE_SI, CDN, nD, nE, SI);
    and (CDN_nD_E_SI, CDN, nD, E, SI);
    and (CDN_D_E_nSI, CDN, D, E, nSI);
    and (CDN_D_nE_nSI, CDN, D, nE, nSI);
    and (CDN_nD_nE_nSI, CDN, nD, nE, nSI);
    and (CDN_D_E_SE, CDN, D, E, SE);
    and (CDN_D_nE_SE, CDN, D, nE, SE);
    and (CDN_nD_nE_SE, CDN, nD, nE, SE);
    and (CDN_nD_E_SE, CDN, nD, E, SE);
    and (D_E_SE_SI, D, E, SE, SI);
    and (D_E_nSE_SI, D, E, nSE, SI);
    and (D_E_nSE_nSI, D, E, nSE, nSI);
    and (nD_E_SE_SI, nD, E, SE, SI);
    and (D_nE_SE_SI, D, nE, SE, SI);
    and (nD_nE_SE_SI, nD, nE, SE, SI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
    and  (D_check, CDN_i, E_d, SE_int_not);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
    and  (D_check, CDN_i, E, SE_int_not);
  `endif
  and  (E_check, CDN_i, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (negedge CDN &&& CP_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_E_SE_SI_SDFCHK, posedge CP &&& D_E_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_E_nSE_SI_SDFCHK, posedge CP &&& D_E_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_E_nSE_nSI_SDFCHK, posedge CP &&& D_E_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_E_SE_SI_SDFCHK, posedge CP &&& nD_E_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nE_SE_SI_SDFCHK, posedge CP &&& D_nE_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_nE_SE_SI_SDFCHK, posedge CP &&& nD_nE_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_E_SE_SI_SDFCHK, posedge CP &&& D_E_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_E_nSE_SI_SDFCHK, posedge CP &&& D_E_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_E_nSE_nSI_SDFCHK, posedge CP &&& D_E_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_E_SE_SI_SDFCHK, posedge CP &&& nD_E_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nE_SE_SI_SDFCHK, posedge CP &&& D_nE_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_nE_SE_SI_SDFCHK, posedge CP &&& nD_nE_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_E_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_E_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_E_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_E_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nE_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_nE_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_E_SE_SI_SDFCHK, posedge CP &&& D_E_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_E_nSE_SI_SDFCHK, posedge CP &&& D_E_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_E_nSE_nSI_SDFCHK, posedge CP &&& D_E_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_E_SE_SI_SDFCHK, posedge CP &&& nD_E_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nE_SE_SI_SDFCHK, posedge CP &&& D_nE_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_nE_SE_SI_SDFCHK, posedge CP &&& nD_nE_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_E_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_E_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_E_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_E_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nE_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_nE_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFCND1 (E, SE, CP, SI, D, CDN, Q, QN);
    input E, SE, CP, SI, D, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire E_d, SE_d, CP_d, SI_d, D_d;
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_E_SE_SI_SDFCHK, CP_D_E_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_E_SE_nSI_SDFCHK, CP_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_E_nSE_SI_SDFCHK, CP_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_E_nSE_nSI_SDFCHK, CP_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_E_SE_SI_SDFCHK, CP_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_E_SE_nSI_SDFCHK, CP_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_E_nSE_SI_SDFCHK, CP_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_E_nSE_nSI_SDFCHK, CP_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nE_SE_SI_SDFCHK, CP_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_nE_SE_nSI_SDFCHK, CP_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nE_nSE_SI_SDFCHK, CP_D_nE_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nE_nSE_nSI_SDFCHK, CP_D_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nE_SE_SI_SDFCHK, CP_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nE_SE_nSI_SDFCHK, CP_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nE_nSE_SI_SDFCHK, CP_nD_nE_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nE_nSE_nSI_SDFCHK, CP_nD_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_E_SE_SI_SDFCHK, nCP_D_E_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_E_SE_nSI_SDFCHK, nCP_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_E_nSE_SI_SDFCHK, nCP_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_E_nSE_nSI_SDFCHK, nCP_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_E_SE_SI_SDFCHK, nCP_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_E_SE_nSI_SDFCHK, nCP_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_E_nSE_SI_SDFCHK, nCP_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_E_nSE_nSI_SDFCHK, nCP_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nE_SE_SI_SDFCHK, nCP_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nE_SE_nSI_SDFCHK, nCP_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nE_nSE_SI_SDFCHK, nCP_D_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nE_nSE_nSI_SDFCHK, nCP_D_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nE_SE_SI_SDFCHK, nCP_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nE_SE_nSI_SDFCHK, nCP_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nE_nSE_SI_SDFCHK, nCP_nD_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nE_nSE_nSI_SDFCHK, nCP_nD_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_E_SE_SI_SDFCHK, CDN_D_E_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_E_nSE_SI_SDFCHK, CDN_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_E_nSE_nSI_SDFCHK, CDN_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_E_SE_SI_SDFCHK, CDN_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nE_SE_SI_SDFCHK, CDN_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SE_SI_SDFCHK, CDN_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_E_SE_nSI_SDFCHK, CDN_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_E_SE_nSI_SDFCHK, CDN_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_E_nSE_SI_SDFCHK, CDN_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_E_nSE_nSI_SDFCHK, CDN_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_nE_SE_nSI_SDFCHK, CDN_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SE_nSI_SDFCHK, CDN_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_E_nSE_SI_SDFCHK, CDN_E_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_E_nSE_nSI_SDFCHK, CDN_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_nE_SI_SDFCHK, CDN_D_nE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SI_SDFCHK, CDN_nD_nE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_E_SI_SDFCHK, CDN_nD_E_SI, 1'b1);
    tsmc_xbuf (CDN_D_E_nSI_SDFCHK, CDN_D_E_nSI, 1'b1);
    tsmc_xbuf (CDN_D_nE_nSI_SDFCHK, CDN_D_nE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nE_nSI_SDFCHK, CDN_nD_nE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_E_SE_SDFCHK, CDN_D_E_SE, 1'b1);
    tsmc_xbuf (CDN_nD_E_SE_SDFCHK, CDN_nD_E_SE, 1'b1);
    tsmc_xbuf (CDN_D_nE_SE_SDFCHK, CDN_D_nE_SE, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SE_SDFCHK, CDN_nD_nE_SE, 1'b1);
    tsmc_xbuf (D_E_SE_SI_SDFCHK, D_E_SE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_SI_SDFCHK, D_E_nSE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_nSI_SDFCHK, D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_E_SE_SI_SDFCHK, nD_E_SE_SI, 1'b1);
    tsmc_xbuf (D_nE_SE_SI_SDFCHK, D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SE_SI_SDFCHK, nD_nE_SE_SI, 1'b1);
  `endif

    not (nE, E);
    not (nSE, SE);
    not (nCP, CP);
    not (nSI, SI);
    not (nD, D);
    and (CP_D_E_SE_SI, CP, D, E, SE, SI);
    and (CP_D_E_SE_nSI, CP, D, E, SE, nSI);
    and (CP_D_E_nSE_SI, CP, D, E, nSE, SI);
    and (CP_D_E_nSE_nSI, CP, D, E, nSE, nSI);
    and (CP_nD_E_SE_SI, CP, nD, E, SE, SI);
    and (CP_nD_E_SE_nSI, CP, nD, E, SE, nSI);
    and (CP_nD_E_nSE_SI, CP, nD, E, nSE, SI);
    and (CP_nD_E_nSE_nSI, CP, nD, E, nSE, nSI);
    and (CP_D_nE_SE_SI, CP, D, nE, SE, SI);
    and (CP_D_nE_SE_nSI, CP, D, nE, SE, nSI);
    and (CP_D_nE_nSE_SI, CP, D, nE, nSE, SI);
    and (CP_D_nE_nSE_nSI, CP, D, nE, nSE, nSI);
    and (CP_nD_nE_SE_SI, CP, nD, nE, SE, SI);
    and (CP_nD_nE_SE_nSI, CP, nD, nE, SE, nSI);
    and (CP_nD_nE_nSE_SI, CP, nD, nE, nSE, SI);
    and (CP_nD_nE_nSE_nSI, CP, nD, nE, nSE, nSI);
    and (nCP_D_E_SE_SI, nCP, D, E, SE, SI);
    and (nCP_D_E_SE_nSI, nCP, D, E, SE, nSI);
    and (nCP_D_E_nSE_SI, nCP, D, E, nSE, SI);
    and (nCP_D_E_nSE_nSI, nCP, D, E, nSE, nSI);
    and (nCP_nD_E_SE_SI, nCP, nD, E, SE, SI);
    and (nCP_nD_E_SE_nSI, nCP, nD, E, SE, nSI);
    and (nCP_nD_E_nSE_SI, nCP, nD, E, nSE, SI);
    and (nCP_nD_E_nSE_nSI, nCP, nD, E, nSE, nSI);
    and (nCP_D_nE_SE_SI, nCP, D, nE, SE, SI);
    and (nCP_D_nE_SE_nSI, nCP, D, nE, SE, nSI);
    and (nCP_D_nE_nSE_SI, nCP, D, nE, nSE, SI);
    and (nCP_D_nE_nSE_nSI, nCP, D, nE, nSE, nSI);
    and (nCP_nD_nE_SE_SI, nCP, nD, nE, SE, SI);
    and (nCP_nD_nE_SE_nSI, nCP, nD, nE, SE, nSI);
    and (nCP_nD_nE_nSE_SI, nCP, nD, nE, nSE, SI);
    and (nCP_nD_nE_nSE_nSI, nCP, nD, nE, nSE, nSI);
    and (CDN_D_E_SE_SI, CDN, D, E, SE, SI);
    and (CDN_D_E_nSE_SI, CDN, D, E, nSE, SI);
    and (CDN_D_E_nSE_nSI, CDN, D, E, nSE, nSI);
    and (CDN_nD_E_SE_SI, CDN, nD, E, SE, SI);
    and (CDN_D_nE_SE_SI, CDN, D, nE, SE, SI);
    and (CDN_nD_nE_SE_SI, CDN, nD, nE, SE, SI);
    and (CDN_D_E_SE_nSI, CDN, D, E, SE, nSI);
    and (CDN_nD_E_SE_nSI, CDN, nD, E, SE, nSI);
    and (CDN_nD_E_nSE_SI, CDN, nD, E, nSE, SI);
    and (CDN_nD_E_nSE_nSI, CDN, nD, E, nSE, nSI);
    and (CDN_D_nE_SE_nSI, CDN, D, nE, SE, nSI);
    and (CDN_nD_nE_SE_nSI, CDN, nD, nE, SE, nSI);
    and (CDN_E_nSE_SI, CDN, E, nSE, SI);
    and (CDN_E_nSE_nSI, CDN, E, nSE, nSI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_D_nE_SI, CDN, D, nE, SI);
    and (CDN_nD_nE_SI, CDN, nD, nE, SI);
    and (CDN_nD_E_SI, CDN, nD, E, SI);
    and (CDN_D_E_nSI, CDN, D, E, nSI);
    and (CDN_D_nE_nSI, CDN, D, nE, nSI);
    and (CDN_nD_nE_nSI, CDN, nD, nE, nSI);
    and (CDN_D_E_SE, CDN, D, E, SE);
    and (CDN_nD_E_SE, CDN, nD, E, SE);
    and (CDN_D_nE_SE, CDN, D, nE, SE);
    and (CDN_nD_nE_SE, CDN, nD, nE, SE);
    and (D_E_SE_SI, D, E, SE, SI);
    and (D_E_nSE_SI, D, E, nSE, SI);
    and (D_E_nSE_nSI, D, E, nSE, nSI);
    and (nD_E_SE_SI, nD, E, SE, SI);
    and (D_nE_SE_SI, D, nE, SE, SI);
    and (nD_nE_SE_SI, nD, nE, SE, SI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
    and  (D_check, CDN_i, E_d, SE_int_not);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
    and  (D_check, CDN_i, E, SE_int_not);
  `endif
  and  (E_check, CDN_i, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (negedge CDN &&& CP_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_E_SE_SI_SDFCHK, posedge CP &&& D_E_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_E_nSE_SI_SDFCHK, posedge CP &&& D_E_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_E_nSE_nSI_SDFCHK, posedge CP &&& D_E_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_E_SE_SI_SDFCHK, posedge CP &&& nD_E_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nE_SE_SI_SDFCHK, posedge CP &&& D_nE_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_nE_SE_SI_SDFCHK, posedge CP &&& nD_nE_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_E_SE_SI_SDFCHK, posedge CP &&& D_E_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_E_nSE_SI_SDFCHK, posedge CP &&& D_E_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_E_nSE_nSI_SDFCHK, posedge CP &&& D_E_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_E_SE_SI_SDFCHK, posedge CP &&& nD_E_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nE_SE_SI_SDFCHK, posedge CP &&& D_nE_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_nE_SE_SI_SDFCHK, posedge CP &&& nD_nE_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_E_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_E_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_E_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_E_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nE_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_nE_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_E_SE_SI_SDFCHK, posedge CP &&& D_E_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_E_nSE_SI_SDFCHK, posedge CP &&& D_E_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_E_nSE_nSI_SDFCHK, posedge CP &&& D_E_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_E_SE_SI_SDFCHK, posedge CP &&& nD_E_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nE_SE_SI_SDFCHK, posedge CP &&& D_nE_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_nE_SE_SI_SDFCHK, posedge CP &&& nD_nE_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_E_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_E_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_E_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_E_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nE_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_nE_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFCND2 (E, SE, CP, SI, D, CDN, Q, QN);
    input E, SE, CP, SI, D, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire E_d, SE_d, CP_d, SI_d, D_d;
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_E_SE_SI_SDFCHK, CP_D_E_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_E_SE_nSI_SDFCHK, CP_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_E_nSE_SI_SDFCHK, CP_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_E_nSE_nSI_SDFCHK, CP_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_E_SE_SI_SDFCHK, CP_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_E_SE_nSI_SDFCHK, CP_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_E_nSE_SI_SDFCHK, CP_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_E_nSE_nSI_SDFCHK, CP_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nE_SE_SI_SDFCHK, CP_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_nE_SE_nSI_SDFCHK, CP_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nE_nSE_SI_SDFCHK, CP_D_nE_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nE_nSE_nSI_SDFCHK, CP_D_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nE_SE_SI_SDFCHK, CP_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nE_SE_nSI_SDFCHK, CP_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nE_nSE_SI_SDFCHK, CP_nD_nE_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nE_nSE_nSI_SDFCHK, CP_nD_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_E_SE_SI_SDFCHK, nCP_D_E_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_E_SE_nSI_SDFCHK, nCP_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_E_nSE_SI_SDFCHK, nCP_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_E_nSE_nSI_SDFCHK, nCP_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_E_SE_SI_SDFCHK, nCP_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_E_SE_nSI_SDFCHK, nCP_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_E_nSE_SI_SDFCHK, nCP_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_E_nSE_nSI_SDFCHK, nCP_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nE_SE_SI_SDFCHK, nCP_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nE_SE_nSI_SDFCHK, nCP_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nE_nSE_SI_SDFCHK, nCP_D_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nE_nSE_nSI_SDFCHK, nCP_D_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nE_SE_SI_SDFCHK, nCP_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nE_SE_nSI_SDFCHK, nCP_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nE_nSE_SI_SDFCHK, nCP_nD_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nE_nSE_nSI_SDFCHK, nCP_nD_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_E_SE_SI_SDFCHK, CDN_D_E_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_E_nSE_SI_SDFCHK, CDN_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_E_nSE_nSI_SDFCHK, CDN_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_E_SE_SI_SDFCHK, CDN_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nE_SE_SI_SDFCHK, CDN_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SE_SI_SDFCHK, CDN_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_E_SE_nSI_SDFCHK, CDN_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_E_SE_nSI_SDFCHK, CDN_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_E_nSE_SI_SDFCHK, CDN_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_E_nSE_nSI_SDFCHK, CDN_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_nE_SE_nSI_SDFCHK, CDN_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SE_nSI_SDFCHK, CDN_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_E_nSE_SI_SDFCHK, CDN_E_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_E_nSE_nSI_SDFCHK, CDN_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_nE_SI_SDFCHK, CDN_D_nE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SI_SDFCHK, CDN_nD_nE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_E_SI_SDFCHK, CDN_nD_E_SI, 1'b1);
    tsmc_xbuf (CDN_D_E_nSI_SDFCHK, CDN_D_E_nSI, 1'b1);
    tsmc_xbuf (CDN_D_nE_nSI_SDFCHK, CDN_D_nE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nE_nSI_SDFCHK, CDN_nD_nE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_E_SE_SDFCHK, CDN_D_E_SE, 1'b1);
    tsmc_xbuf (CDN_nD_E_SE_SDFCHK, CDN_nD_E_SE, 1'b1);
    tsmc_xbuf (CDN_D_nE_SE_SDFCHK, CDN_D_nE_SE, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SE_SDFCHK, CDN_nD_nE_SE, 1'b1);
    tsmc_xbuf (D_E_SE_SI_SDFCHK, D_E_SE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_SI_SDFCHK, D_E_nSE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_nSI_SDFCHK, D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_E_SE_SI_SDFCHK, nD_E_SE_SI, 1'b1);
    tsmc_xbuf (D_nE_SE_SI_SDFCHK, D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SE_SI_SDFCHK, nD_nE_SE_SI, 1'b1);
  `endif

    not (nE, E);
    not (nSE, SE);
    not (nCP, CP);
    not (nSI, SI);
    not (nD, D);
    and (CP_D_E_SE_SI, CP, D, E, SE, SI);
    and (CP_D_E_SE_nSI, CP, D, E, SE, nSI);
    and (CP_D_E_nSE_SI, CP, D, E, nSE, SI);
    and (CP_D_E_nSE_nSI, CP, D, E, nSE, nSI);
    and (CP_nD_E_SE_SI, CP, nD, E, SE, SI);
    and (CP_nD_E_SE_nSI, CP, nD, E, SE, nSI);
    and (CP_nD_E_nSE_SI, CP, nD, E, nSE, SI);
    and (CP_nD_E_nSE_nSI, CP, nD, E, nSE, nSI);
    and (CP_D_nE_SE_SI, CP, D, nE, SE, SI);
    and (CP_D_nE_SE_nSI, CP, D, nE, SE, nSI);
    and (CP_D_nE_nSE_SI, CP, D, nE, nSE, SI);
    and (CP_D_nE_nSE_nSI, CP, D, nE, nSE, nSI);
    and (CP_nD_nE_SE_SI, CP, nD, nE, SE, SI);
    and (CP_nD_nE_SE_nSI, CP, nD, nE, SE, nSI);
    and (CP_nD_nE_nSE_SI, CP, nD, nE, nSE, SI);
    and (CP_nD_nE_nSE_nSI, CP, nD, nE, nSE, nSI);
    and (nCP_D_E_SE_SI, nCP, D, E, SE, SI);
    and (nCP_D_E_SE_nSI, nCP, D, E, SE, nSI);
    and (nCP_D_E_nSE_SI, nCP, D, E, nSE, SI);
    and (nCP_D_E_nSE_nSI, nCP, D, E, nSE, nSI);
    and (nCP_nD_E_SE_SI, nCP, nD, E, SE, SI);
    and (nCP_nD_E_SE_nSI, nCP, nD, E, SE, nSI);
    and (nCP_nD_E_nSE_SI, nCP, nD, E, nSE, SI);
    and (nCP_nD_E_nSE_nSI, nCP, nD, E, nSE, nSI);
    and (nCP_D_nE_SE_SI, nCP, D, nE, SE, SI);
    and (nCP_D_nE_SE_nSI, nCP, D, nE, SE, nSI);
    and (nCP_D_nE_nSE_SI, nCP, D, nE, nSE, SI);
    and (nCP_D_nE_nSE_nSI, nCP, D, nE, nSE, nSI);
    and (nCP_nD_nE_SE_SI, nCP, nD, nE, SE, SI);
    and (nCP_nD_nE_SE_nSI, nCP, nD, nE, SE, nSI);
    and (nCP_nD_nE_nSE_SI, nCP, nD, nE, nSE, SI);
    and (nCP_nD_nE_nSE_nSI, nCP, nD, nE, nSE, nSI);
    and (CDN_D_E_SE_SI, CDN, D, E, SE, SI);
    and (CDN_D_E_nSE_SI, CDN, D, E, nSE, SI);
    and (CDN_D_E_nSE_nSI, CDN, D, E, nSE, nSI);
    and (CDN_nD_E_SE_SI, CDN, nD, E, SE, SI);
    and (CDN_D_nE_SE_SI, CDN, D, nE, SE, SI);
    and (CDN_nD_nE_SE_SI, CDN, nD, nE, SE, SI);
    and (CDN_D_E_SE_nSI, CDN, D, E, SE, nSI);
    and (CDN_nD_E_SE_nSI, CDN, nD, E, SE, nSI);
    and (CDN_nD_E_nSE_SI, CDN, nD, E, nSE, SI);
    and (CDN_nD_E_nSE_nSI, CDN, nD, E, nSE, nSI);
    and (CDN_D_nE_SE_nSI, CDN, D, nE, SE, nSI);
    and (CDN_nD_nE_SE_nSI, CDN, nD, nE, SE, nSI);
    and (CDN_E_nSE_SI, CDN, E, nSE, SI);
    and (CDN_E_nSE_nSI, CDN, E, nSE, nSI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_D_nE_SI, CDN, D, nE, SI);
    and (CDN_nD_nE_SI, CDN, nD, nE, SI);
    and (CDN_nD_E_SI, CDN, nD, E, SI);
    and (CDN_D_E_nSI, CDN, D, E, nSI);
    and (CDN_D_nE_nSI, CDN, D, nE, nSI);
    and (CDN_nD_nE_nSI, CDN, nD, nE, nSI);
    and (CDN_D_E_SE, CDN, D, E, SE);
    and (CDN_nD_E_SE, CDN, nD, E, SE);
    and (CDN_D_nE_SE, CDN, D, nE, SE);
    and (CDN_nD_nE_SE, CDN, nD, nE, SE);
    and (D_E_SE_SI, D, E, SE, SI);
    and (D_E_nSE_SI, D, E, nSE, SI);
    and (D_E_nSE_nSI, D, E, nSE, nSI);
    and (nD_E_SE_SI, nD, E, SE, SI);
    and (D_nE_SE_SI, D, nE, SE, SI);
    and (nD_nE_SE_SI, nD, nE, SE, SI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
    and  (D_check, CDN_i, E_d, SE_int_not);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
    and  (D_check, CDN_i, E, SE_int_not);
  `endif
  and  (E_check, CDN_i, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (negedge CDN &&& CP_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_E_SE_SI_SDFCHK, posedge CP &&& D_E_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_E_nSE_SI_SDFCHK, posedge CP &&& D_E_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_E_nSE_nSI_SDFCHK, posedge CP &&& D_E_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_E_SE_SI_SDFCHK, posedge CP &&& nD_E_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nE_SE_SI_SDFCHK, posedge CP &&& D_nE_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_nE_SE_SI_SDFCHK, posedge CP &&& nD_nE_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_E_SE_SI_SDFCHK, posedge CP &&& D_E_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_E_nSE_SI_SDFCHK, posedge CP &&& D_E_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_E_nSE_nSI_SDFCHK, posedge CP &&& D_E_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_E_SE_SI_SDFCHK, posedge CP &&& nD_E_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nE_SE_SI_SDFCHK, posedge CP &&& D_nE_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_nE_SE_SI_SDFCHK, posedge CP &&& nD_nE_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_E_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_E_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_E_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_E_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nE_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_nE_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_E_SE_SI_SDFCHK, posedge CP &&& D_E_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_E_nSE_SI_SDFCHK, posedge CP &&& D_E_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_E_nSE_nSI_SDFCHK, posedge CP &&& D_E_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_E_SE_SI_SDFCHK, posedge CP &&& nD_E_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nE_SE_SI_SDFCHK, posedge CP &&& D_nE_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_nE_SE_SI_SDFCHK, posedge CP &&& nD_nE_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_E_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_E_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_E_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_E_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nE_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_nE_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFCND4 (E, SE, CP, SI, D, CDN, Q, QN);
    input E, SE, CP, SI, D, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire E_d, SE_d, CP_d, SI_d, D_d;
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_E_SE_SI_SDFCHK, CP_D_E_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_E_SE_nSI_SDFCHK, CP_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_E_nSE_SI_SDFCHK, CP_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_E_nSE_nSI_SDFCHK, CP_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_E_SE_SI_SDFCHK, CP_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_E_SE_nSI_SDFCHK, CP_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_E_nSE_SI_SDFCHK, CP_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_E_nSE_nSI_SDFCHK, CP_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nE_SE_SI_SDFCHK, CP_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_nE_SE_nSI_SDFCHK, CP_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nE_nSE_SI_SDFCHK, CP_D_nE_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nE_nSE_nSI_SDFCHK, CP_D_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nE_SE_SI_SDFCHK, CP_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nE_SE_nSI_SDFCHK, CP_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nE_nSE_SI_SDFCHK, CP_nD_nE_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nE_nSE_nSI_SDFCHK, CP_nD_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_E_SE_SI_SDFCHK, nCP_D_E_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_E_SE_nSI_SDFCHK, nCP_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_E_nSE_SI_SDFCHK, nCP_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_E_nSE_nSI_SDFCHK, nCP_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_E_SE_SI_SDFCHK, nCP_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_E_SE_nSI_SDFCHK, nCP_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_E_nSE_SI_SDFCHK, nCP_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_E_nSE_nSI_SDFCHK, nCP_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nE_SE_SI_SDFCHK, nCP_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nE_SE_nSI_SDFCHK, nCP_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nE_nSE_SI_SDFCHK, nCP_D_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nE_nSE_nSI_SDFCHK, nCP_D_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nE_SE_SI_SDFCHK, nCP_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nE_SE_nSI_SDFCHK, nCP_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nE_nSE_SI_SDFCHK, nCP_nD_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nE_nSE_nSI_SDFCHK, nCP_nD_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_E_SE_SI_SDFCHK, CDN_D_E_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_E_nSE_SI_SDFCHK, CDN_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_E_nSE_nSI_SDFCHK, CDN_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_E_SE_SI_SDFCHK, CDN_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nE_SE_SI_SDFCHK, CDN_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SE_SI_SDFCHK, CDN_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_E_SE_nSI_SDFCHK, CDN_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_E_SE_nSI_SDFCHK, CDN_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_E_nSE_SI_SDFCHK, CDN_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_E_nSE_nSI_SDFCHK, CDN_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_nE_SE_nSI_SDFCHK, CDN_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SE_nSI_SDFCHK, CDN_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_E_nSE_SI_SDFCHK, CDN_E_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_E_nSE_nSI_SDFCHK, CDN_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_nE_SI_SDFCHK, CDN_D_nE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SI_SDFCHK, CDN_nD_nE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_E_SI_SDFCHK, CDN_nD_E_SI, 1'b1);
    tsmc_xbuf (CDN_D_E_nSI_SDFCHK, CDN_D_E_nSI, 1'b1);
    tsmc_xbuf (CDN_D_nE_nSI_SDFCHK, CDN_D_nE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nE_nSI_SDFCHK, CDN_nD_nE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_E_SE_SDFCHK, CDN_D_E_SE, 1'b1);
    tsmc_xbuf (CDN_nD_E_SE_SDFCHK, CDN_nD_E_SE, 1'b1);
    tsmc_xbuf (CDN_D_nE_SE_SDFCHK, CDN_D_nE_SE, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SE_SDFCHK, CDN_nD_nE_SE, 1'b1);
    tsmc_xbuf (D_E_SE_SI_SDFCHK, D_E_SE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_SI_SDFCHK, D_E_nSE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_nSI_SDFCHK, D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_E_SE_SI_SDFCHK, nD_E_SE_SI, 1'b1);
    tsmc_xbuf (D_nE_SE_SI_SDFCHK, D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SE_SI_SDFCHK, nD_nE_SE_SI, 1'b1);
  `endif

    not (nE, E);
    not (nSE, SE);
    not (nCP, CP);
    not (nSI, SI);
    not (nD, D);
    and (CP_D_E_SE_SI, CP, D, E, SE, SI);
    and (CP_D_E_SE_nSI, CP, D, E, SE, nSI);
    and (CP_D_E_nSE_SI, CP, D, E, nSE, SI);
    and (CP_D_E_nSE_nSI, CP, D, E, nSE, nSI);
    and (CP_nD_E_SE_SI, CP, nD, E, SE, SI);
    and (CP_nD_E_SE_nSI, CP, nD, E, SE, nSI);
    and (CP_nD_E_nSE_SI, CP, nD, E, nSE, SI);
    and (CP_nD_E_nSE_nSI, CP, nD, E, nSE, nSI);
    and (CP_D_nE_SE_SI, CP, D, nE, SE, SI);
    and (CP_D_nE_SE_nSI, CP, D, nE, SE, nSI);
    and (CP_D_nE_nSE_SI, CP, D, nE, nSE, SI);
    and (CP_D_nE_nSE_nSI, CP, D, nE, nSE, nSI);
    and (CP_nD_nE_SE_SI, CP, nD, nE, SE, SI);
    and (CP_nD_nE_SE_nSI, CP, nD, nE, SE, nSI);
    and (CP_nD_nE_nSE_SI, CP, nD, nE, nSE, SI);
    and (CP_nD_nE_nSE_nSI, CP, nD, nE, nSE, nSI);
    and (nCP_D_E_SE_SI, nCP, D, E, SE, SI);
    and (nCP_D_E_SE_nSI, nCP, D, E, SE, nSI);
    and (nCP_D_E_nSE_SI, nCP, D, E, nSE, SI);
    and (nCP_D_E_nSE_nSI, nCP, D, E, nSE, nSI);
    and (nCP_nD_E_SE_SI, nCP, nD, E, SE, SI);
    and (nCP_nD_E_SE_nSI, nCP, nD, E, SE, nSI);
    and (nCP_nD_E_nSE_SI, nCP, nD, E, nSE, SI);
    and (nCP_nD_E_nSE_nSI, nCP, nD, E, nSE, nSI);
    and (nCP_D_nE_SE_SI, nCP, D, nE, SE, SI);
    and (nCP_D_nE_SE_nSI, nCP, D, nE, SE, nSI);
    and (nCP_D_nE_nSE_SI, nCP, D, nE, nSE, SI);
    and (nCP_D_nE_nSE_nSI, nCP, D, nE, nSE, nSI);
    and (nCP_nD_nE_SE_SI, nCP, nD, nE, SE, SI);
    and (nCP_nD_nE_SE_nSI, nCP, nD, nE, SE, nSI);
    and (nCP_nD_nE_nSE_SI, nCP, nD, nE, nSE, SI);
    and (nCP_nD_nE_nSE_nSI, nCP, nD, nE, nSE, nSI);
    and (CDN_D_E_SE_SI, CDN, D, E, SE, SI);
    and (CDN_D_E_nSE_SI, CDN, D, E, nSE, SI);
    and (CDN_D_E_nSE_nSI, CDN, D, E, nSE, nSI);
    and (CDN_nD_E_SE_SI, CDN, nD, E, SE, SI);
    and (CDN_D_nE_SE_SI, CDN, D, nE, SE, SI);
    and (CDN_nD_nE_SE_SI, CDN, nD, nE, SE, SI);
    and (CDN_D_E_SE_nSI, CDN, D, E, SE, nSI);
    and (CDN_nD_E_SE_nSI, CDN, nD, E, SE, nSI);
    and (CDN_nD_E_nSE_SI, CDN, nD, E, nSE, SI);
    and (CDN_nD_E_nSE_nSI, CDN, nD, E, nSE, nSI);
    and (CDN_D_nE_SE_nSI, CDN, D, nE, SE, nSI);
    and (CDN_nD_nE_SE_nSI, CDN, nD, nE, SE, nSI);
    and (CDN_E_nSE_SI, CDN, E, nSE, SI);
    and (CDN_E_nSE_nSI, CDN, E, nSE, nSI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_D_nE_SI, CDN, D, nE, SI);
    and (CDN_nD_nE_SI, CDN, nD, nE, SI);
    and (CDN_nD_E_SI, CDN, nD, E, SI);
    and (CDN_D_E_nSI, CDN, D, E, nSI);
    and (CDN_D_nE_nSI, CDN, D, nE, nSI);
    and (CDN_nD_nE_nSI, CDN, nD, nE, nSI);
    and (CDN_D_E_SE, CDN, D, E, SE);
    and (CDN_nD_E_SE, CDN, nD, E, SE);
    and (CDN_D_nE_SE, CDN, D, nE, SE);
    and (CDN_nD_nE_SE, CDN, nD, nE, SE);
    and (D_E_SE_SI, D, E, SE, SI);
    and (D_E_nSE_SI, D, E, nSE, SI);
    and (D_E_nSE_nSI, D, E, nSE, nSI);
    and (nD_E_SE_SI, nD, E, SE, SI);
    and (D_nE_SE_SI, D, nE, SE, SI);
    and (nD_nE_SE_SI, nD, nE, SE, SI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
    and  (D_check, CDN_i, E_d, SE_int_not);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
    and  (D_check, CDN_i, E, SE_int_not);
  `endif
  and  (E_check, CDN_i, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (negedge CDN &&& CP_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_E_SE_SI_SDFCHK, posedge CP &&& D_E_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_E_nSE_SI_SDFCHK, posedge CP &&& D_E_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_E_nSE_nSI_SDFCHK, posedge CP &&& D_E_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_E_SE_SI_SDFCHK, posedge CP &&& nD_E_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nE_SE_SI_SDFCHK, posedge CP &&& D_nE_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_nE_SE_SI_SDFCHK, posedge CP &&& nD_nE_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_E_SE_SI_SDFCHK, posedge CP &&& D_E_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_E_nSE_SI_SDFCHK, posedge CP &&& D_E_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_E_nSE_nSI_SDFCHK, posedge CP &&& D_E_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_E_SE_SI_SDFCHK, posedge CP &&& nD_E_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nE_SE_SI_SDFCHK, posedge CP &&& D_nE_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_nE_SE_SI_SDFCHK, posedge CP &&& nD_nE_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_E_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_E_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_E_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_E_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nE_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_nE_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_E_SE_SI_SDFCHK, posedge CP &&& D_E_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_E_nSE_SI_SDFCHK, posedge CP &&& D_E_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_E_nSE_nSI_SDFCHK, posedge CP &&& D_E_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_E_SE_SI_SDFCHK, posedge CP &&& nD_E_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nE_SE_SI_SDFCHK, posedge CP &&& D_nE_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_nE_SE_SI_SDFCHK, posedge CP &&& nD_nE_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_E_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_E_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_E_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_E_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nE_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_nE_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFCNQD0 (E, SE, CP, SI, D, CDN, Q);
    input E, SE, CP, SI, D, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire E_d, SE_d, CP_d, SI_d, D_d;
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_E_SE_SI_SDFCHK, CP_D_E_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_E_SE_nSI_SDFCHK, CP_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_E_nSE_SI_SDFCHK, CP_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_E_nSE_nSI_SDFCHK, CP_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_E_SE_SI_SDFCHK, CP_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_E_SE_nSI_SDFCHK, CP_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_E_nSE_SI_SDFCHK, CP_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_E_nSE_nSI_SDFCHK, CP_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nE_SE_SI_SDFCHK, CP_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_nE_SE_nSI_SDFCHK, CP_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nE_nSE_SI_SDFCHK, CP_D_nE_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nE_nSE_nSI_SDFCHK, CP_D_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nE_SE_SI_SDFCHK, CP_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nE_SE_nSI_SDFCHK, CP_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nE_nSE_SI_SDFCHK, CP_nD_nE_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nE_nSE_nSI_SDFCHK, CP_nD_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_E_SE_SI_SDFCHK, nCP_D_E_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_E_SE_nSI_SDFCHK, nCP_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_E_nSE_SI_SDFCHK, nCP_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_E_nSE_nSI_SDFCHK, nCP_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_E_SE_SI_SDFCHK, nCP_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_E_SE_nSI_SDFCHK, nCP_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_E_nSE_SI_SDFCHK, nCP_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_E_nSE_nSI_SDFCHK, nCP_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nE_SE_SI_SDFCHK, nCP_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nE_SE_nSI_SDFCHK, nCP_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nE_nSE_SI_SDFCHK, nCP_D_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nE_nSE_nSI_SDFCHK, nCP_D_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nE_SE_SI_SDFCHK, nCP_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nE_SE_nSI_SDFCHK, nCP_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nE_nSE_SI_SDFCHK, nCP_nD_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nE_nSE_nSI_SDFCHK, nCP_nD_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_E_SE_SI_SDFCHK, CDN_D_E_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_E_nSE_SI_SDFCHK, CDN_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_E_nSE_nSI_SDFCHK, CDN_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_E_SE_SI_SDFCHK, CDN_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nE_SE_SI_SDFCHK, CDN_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SE_SI_SDFCHK, CDN_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_E_SE_nSI_SDFCHK, CDN_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_E_SE_nSI_SDFCHK, CDN_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_E_nSE_SI_SDFCHK, CDN_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_E_nSE_nSI_SDFCHK, CDN_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_nE_SE_nSI_SDFCHK, CDN_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SE_nSI_SDFCHK, CDN_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_E_nSE_SI_SDFCHK, CDN_E_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_E_nSE_nSI_SDFCHK, CDN_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_nE_SI_SDFCHK, CDN_D_nE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SI_SDFCHK, CDN_nD_nE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_E_SI_SDFCHK, CDN_nD_E_SI, 1'b1);
    tsmc_xbuf (CDN_D_E_nSI_SDFCHK, CDN_D_E_nSI, 1'b1);
    tsmc_xbuf (CDN_D_nE_nSI_SDFCHK, CDN_D_nE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nE_nSI_SDFCHK, CDN_nD_nE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_E_SE_SDFCHK, CDN_D_E_SE, 1'b1);
    tsmc_xbuf (CDN_D_nE_SE_SDFCHK, CDN_D_nE_SE, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SE_SDFCHK, CDN_nD_nE_SE, 1'b1);
    tsmc_xbuf (CDN_nD_E_SE_SDFCHK, CDN_nD_E_SE, 1'b1);
    tsmc_xbuf (D_E_SE_SI_SDFCHK, D_E_SE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_SI_SDFCHK, D_E_nSE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_nSI_SDFCHK, D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_E_SE_SI_SDFCHK, nD_E_SE_SI, 1'b1);
    tsmc_xbuf (D_nE_SE_SI_SDFCHK, D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SE_SI_SDFCHK, nD_nE_SE_SI, 1'b1);
  `endif

    not (nE, E);
    not (nSE, SE);
    not (nCP, CP);
    not (nSI, SI);
    not (nD, D);
    and (CP_D_E_SE_SI, CP, D, E, SE, SI);
    and (CP_D_E_SE_nSI, CP, D, E, SE, nSI);
    and (CP_D_E_nSE_SI, CP, D, E, nSE, SI);
    and (CP_D_E_nSE_nSI, CP, D, E, nSE, nSI);
    and (CP_nD_E_SE_SI, CP, nD, E, SE, SI);
    and (CP_nD_E_SE_nSI, CP, nD, E, SE, nSI);
    and (CP_nD_E_nSE_SI, CP, nD, E, nSE, SI);
    and (CP_nD_E_nSE_nSI, CP, nD, E, nSE, nSI);
    and (CP_D_nE_SE_SI, CP, D, nE, SE, SI);
    and (CP_D_nE_SE_nSI, CP, D, nE, SE, nSI);
    and (CP_D_nE_nSE_SI, CP, D, nE, nSE, SI);
    and (CP_D_nE_nSE_nSI, CP, D, nE, nSE, nSI);
    and (CP_nD_nE_SE_SI, CP, nD, nE, SE, SI);
    and (CP_nD_nE_SE_nSI, CP, nD, nE, SE, nSI);
    and (CP_nD_nE_nSE_SI, CP, nD, nE, nSE, SI);
    and (CP_nD_nE_nSE_nSI, CP, nD, nE, nSE, nSI);
    and (nCP_D_E_SE_SI, nCP, D, E, SE, SI);
    and (nCP_D_E_SE_nSI, nCP, D, E, SE, nSI);
    and (nCP_D_E_nSE_SI, nCP, D, E, nSE, SI);
    and (nCP_D_E_nSE_nSI, nCP, D, E, nSE, nSI);
    and (nCP_nD_E_SE_SI, nCP, nD, E, SE, SI);
    and (nCP_nD_E_SE_nSI, nCP, nD, E, SE, nSI);
    and (nCP_nD_E_nSE_SI, nCP, nD, E, nSE, SI);
    and (nCP_nD_E_nSE_nSI, nCP, nD, E, nSE, nSI);
    and (nCP_D_nE_SE_SI, nCP, D, nE, SE, SI);
    and (nCP_D_nE_SE_nSI, nCP, D, nE, SE, nSI);
    and (nCP_D_nE_nSE_SI, nCP, D, nE, nSE, SI);
    and (nCP_D_nE_nSE_nSI, nCP, D, nE, nSE, nSI);
    and (nCP_nD_nE_SE_SI, nCP, nD, nE, SE, SI);
    and (nCP_nD_nE_SE_nSI, nCP, nD, nE, SE, nSI);
    and (nCP_nD_nE_nSE_SI, nCP, nD, nE, nSE, SI);
    and (nCP_nD_nE_nSE_nSI, nCP, nD, nE, nSE, nSI);
    and (CDN_D_E_SE_SI, CDN, D, E, SE, SI);
    and (CDN_D_E_nSE_SI, CDN, D, E, nSE, SI);
    and (CDN_D_E_nSE_nSI, CDN, D, E, nSE, nSI);
    and (CDN_nD_E_SE_SI, CDN, nD, E, SE, SI);
    and (CDN_D_nE_SE_SI, CDN, D, nE, SE, SI);
    and (CDN_nD_nE_SE_SI, CDN, nD, nE, SE, SI);
    and (CDN_D_E_SE_nSI, CDN, D, E, SE, nSI);
    and (CDN_nD_E_SE_nSI, CDN, nD, E, SE, nSI);
    and (CDN_nD_E_nSE_SI, CDN, nD, E, nSE, SI);
    and (CDN_nD_E_nSE_nSI, CDN, nD, E, nSE, nSI);
    and (CDN_D_nE_SE_nSI, CDN, D, nE, SE, nSI);
    and (CDN_nD_nE_SE_nSI, CDN, nD, nE, SE, nSI);
    and (CDN_E_nSE_SI, CDN, E, nSE, SI);
    and (CDN_E_nSE_nSI, CDN, E, nSE, nSI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_D_nE_SI, CDN, D, nE, SI);
    and (CDN_nD_nE_SI, CDN, nD, nE, SI);
    and (CDN_nD_E_SI, CDN, nD, E, SI);
    and (CDN_D_E_nSI, CDN, D, E, nSI);
    and (CDN_D_nE_nSI, CDN, D, nE, nSI);
    and (CDN_nD_nE_nSI, CDN, nD, nE, nSI);
    and (CDN_D_E_SE, CDN, D, E, SE);
    and (CDN_D_nE_SE, CDN, D, nE, SE);
    and (CDN_nD_nE_SE, CDN, nD, nE, SE);
    and (CDN_nD_E_SE, CDN, nD, E, SE);
    and (D_E_SE_SI, D, E, SE, SI);
    and (D_E_nSE_SI, D, E, nSE, SI);
    and (D_E_nSE_nSI, D, E, nSE, nSI);
    and (nD_E_SE_SI, nD, E, SE, SI);
    and (D_nE_SE_SI, D, nE, SE, SI);
    and (nD_nE_SE_SI, nD, nE, SE, SI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
    and  (D_check, CDN_i, E_d, SE_int_not);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
    and  (D_check, CDN_i, E, SE_int_not);
  `endif
  and  (E_check, CDN_i, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (negedge CDN &&& CP_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_E_SE_SI_SDFCHK, posedge CP &&& D_E_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_E_nSE_SI_SDFCHK, posedge CP &&& D_E_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_E_nSE_nSI_SDFCHK, posedge CP &&& D_E_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_E_SE_SI_SDFCHK, posedge CP &&& nD_E_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nE_SE_SI_SDFCHK, posedge CP &&& D_nE_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_nE_SE_SI_SDFCHK, posedge CP &&& nD_nE_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_E_SE_SI_SDFCHK, posedge CP &&& D_E_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_E_nSE_SI_SDFCHK, posedge CP &&& D_E_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_E_nSE_nSI_SDFCHK, posedge CP &&& D_E_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_E_SE_SI_SDFCHK, posedge CP &&& nD_E_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nE_SE_SI_SDFCHK, posedge CP &&& D_nE_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_nE_SE_SI_SDFCHK, posedge CP &&& nD_nE_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_E_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_E_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_E_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_E_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nE_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_nE_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_E_SE_SI_SDFCHK, posedge CP &&& D_E_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_E_nSE_SI_SDFCHK, posedge CP &&& D_E_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_E_nSE_nSI_SDFCHK, posedge CP &&& D_E_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_E_SE_SI_SDFCHK, posedge CP &&& nD_E_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nE_SE_SI_SDFCHK, posedge CP &&& D_nE_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_nE_SE_SI_SDFCHK, posedge CP &&& nD_nE_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_E_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_E_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_E_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_E_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nE_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_nE_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFCNQD1 (E, SE, CP, SI, D, CDN, Q);
    input E, SE, CP, SI, D, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire E_d, SE_d, CP_d, SI_d, D_d;
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_E_SE_SI_SDFCHK, CP_D_E_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_E_SE_nSI_SDFCHK, CP_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_E_nSE_SI_SDFCHK, CP_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_E_nSE_nSI_SDFCHK, CP_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_E_SE_SI_SDFCHK, CP_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_E_SE_nSI_SDFCHK, CP_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_E_nSE_SI_SDFCHK, CP_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_E_nSE_nSI_SDFCHK, CP_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nE_SE_SI_SDFCHK, CP_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_nE_SE_nSI_SDFCHK, CP_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nE_nSE_SI_SDFCHK, CP_D_nE_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nE_nSE_nSI_SDFCHK, CP_D_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nE_SE_SI_SDFCHK, CP_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nE_SE_nSI_SDFCHK, CP_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nE_nSE_SI_SDFCHK, CP_nD_nE_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nE_nSE_nSI_SDFCHK, CP_nD_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_E_SE_SI_SDFCHK, nCP_D_E_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_E_SE_nSI_SDFCHK, nCP_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_E_nSE_SI_SDFCHK, nCP_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_E_nSE_nSI_SDFCHK, nCP_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_E_SE_SI_SDFCHK, nCP_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_E_SE_nSI_SDFCHK, nCP_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_E_nSE_SI_SDFCHK, nCP_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_E_nSE_nSI_SDFCHK, nCP_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nE_SE_SI_SDFCHK, nCP_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nE_SE_nSI_SDFCHK, nCP_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nE_nSE_SI_SDFCHK, nCP_D_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nE_nSE_nSI_SDFCHK, nCP_D_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nE_SE_SI_SDFCHK, nCP_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nE_SE_nSI_SDFCHK, nCP_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nE_nSE_SI_SDFCHK, nCP_nD_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nE_nSE_nSI_SDFCHK, nCP_nD_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_E_SE_SI_SDFCHK, CDN_D_E_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_E_nSE_SI_SDFCHK, CDN_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_E_nSE_nSI_SDFCHK, CDN_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_E_SE_SI_SDFCHK, CDN_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nE_SE_SI_SDFCHK, CDN_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SE_SI_SDFCHK, CDN_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_E_SE_nSI_SDFCHK, CDN_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_E_SE_nSI_SDFCHK, CDN_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_E_nSE_SI_SDFCHK, CDN_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_E_nSE_nSI_SDFCHK, CDN_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_nE_SE_nSI_SDFCHK, CDN_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SE_nSI_SDFCHK, CDN_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_E_nSE_SI_SDFCHK, CDN_E_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_E_nSE_nSI_SDFCHK, CDN_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_nE_SI_SDFCHK, CDN_D_nE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SI_SDFCHK, CDN_nD_nE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_E_SI_SDFCHK, CDN_nD_E_SI, 1'b1);
    tsmc_xbuf (CDN_D_E_nSI_SDFCHK, CDN_D_E_nSI, 1'b1);
    tsmc_xbuf (CDN_D_nE_nSI_SDFCHK, CDN_D_nE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nE_nSI_SDFCHK, CDN_nD_nE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_E_SE_SDFCHK, CDN_D_E_SE, 1'b1);
    tsmc_xbuf (CDN_nD_E_SE_SDFCHK, CDN_nD_E_SE, 1'b1);
    tsmc_xbuf (CDN_D_nE_SE_SDFCHK, CDN_D_nE_SE, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SE_SDFCHK, CDN_nD_nE_SE, 1'b1);
    tsmc_xbuf (D_E_SE_SI_SDFCHK, D_E_SE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_SI_SDFCHK, D_E_nSE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_nSI_SDFCHK, D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_E_SE_SI_SDFCHK, nD_E_SE_SI, 1'b1);
    tsmc_xbuf (D_nE_SE_SI_SDFCHK, D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SE_SI_SDFCHK, nD_nE_SE_SI, 1'b1);
  `endif

    not (nE, E);
    not (nSE, SE);
    not (nCP, CP);
    not (nSI, SI);
    not (nD, D);
    and (CP_D_E_SE_SI, CP, D, E, SE, SI);
    and (CP_D_E_SE_nSI, CP, D, E, SE, nSI);
    and (CP_D_E_nSE_SI, CP, D, E, nSE, SI);
    and (CP_D_E_nSE_nSI, CP, D, E, nSE, nSI);
    and (CP_nD_E_SE_SI, CP, nD, E, SE, SI);
    and (CP_nD_E_SE_nSI, CP, nD, E, SE, nSI);
    and (CP_nD_E_nSE_SI, CP, nD, E, nSE, SI);
    and (CP_nD_E_nSE_nSI, CP, nD, E, nSE, nSI);
    and (CP_D_nE_SE_SI, CP, D, nE, SE, SI);
    and (CP_D_nE_SE_nSI, CP, D, nE, SE, nSI);
    and (CP_D_nE_nSE_SI, CP, D, nE, nSE, SI);
    and (CP_D_nE_nSE_nSI, CP, D, nE, nSE, nSI);
    and (CP_nD_nE_SE_SI, CP, nD, nE, SE, SI);
    and (CP_nD_nE_SE_nSI, CP, nD, nE, SE, nSI);
    and (CP_nD_nE_nSE_SI, CP, nD, nE, nSE, SI);
    and (CP_nD_nE_nSE_nSI, CP, nD, nE, nSE, nSI);
    and (nCP_D_E_SE_SI, nCP, D, E, SE, SI);
    and (nCP_D_E_SE_nSI, nCP, D, E, SE, nSI);
    and (nCP_D_E_nSE_SI, nCP, D, E, nSE, SI);
    and (nCP_D_E_nSE_nSI, nCP, D, E, nSE, nSI);
    and (nCP_nD_E_SE_SI, nCP, nD, E, SE, SI);
    and (nCP_nD_E_SE_nSI, nCP, nD, E, SE, nSI);
    and (nCP_nD_E_nSE_SI, nCP, nD, E, nSE, SI);
    and (nCP_nD_E_nSE_nSI, nCP, nD, E, nSE, nSI);
    and (nCP_D_nE_SE_SI, nCP, D, nE, SE, SI);
    and (nCP_D_nE_SE_nSI, nCP, D, nE, SE, nSI);
    and (nCP_D_nE_nSE_SI, nCP, D, nE, nSE, SI);
    and (nCP_D_nE_nSE_nSI, nCP, D, nE, nSE, nSI);
    and (nCP_nD_nE_SE_SI, nCP, nD, nE, SE, SI);
    and (nCP_nD_nE_SE_nSI, nCP, nD, nE, SE, nSI);
    and (nCP_nD_nE_nSE_SI, nCP, nD, nE, nSE, SI);
    and (nCP_nD_nE_nSE_nSI, nCP, nD, nE, nSE, nSI);
    and (CDN_D_E_SE_SI, CDN, D, E, SE, SI);
    and (CDN_D_E_nSE_SI, CDN, D, E, nSE, SI);
    and (CDN_D_E_nSE_nSI, CDN, D, E, nSE, nSI);
    and (CDN_nD_E_SE_SI, CDN, nD, E, SE, SI);
    and (CDN_D_nE_SE_SI, CDN, D, nE, SE, SI);
    and (CDN_nD_nE_SE_SI, CDN, nD, nE, SE, SI);
    and (CDN_D_E_SE_nSI, CDN, D, E, SE, nSI);
    and (CDN_nD_E_SE_nSI, CDN, nD, E, SE, nSI);
    and (CDN_nD_E_nSE_SI, CDN, nD, E, nSE, SI);
    and (CDN_nD_E_nSE_nSI, CDN, nD, E, nSE, nSI);
    and (CDN_D_nE_SE_nSI, CDN, D, nE, SE, nSI);
    and (CDN_nD_nE_SE_nSI, CDN, nD, nE, SE, nSI);
    and (CDN_E_nSE_SI, CDN, E, nSE, SI);
    and (CDN_E_nSE_nSI, CDN, E, nSE, nSI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_D_nE_SI, CDN, D, nE, SI);
    and (CDN_nD_nE_SI, CDN, nD, nE, SI);
    and (CDN_nD_E_SI, CDN, nD, E, SI);
    and (CDN_D_E_nSI, CDN, D, E, nSI);
    and (CDN_D_nE_nSI, CDN, D, nE, nSI);
    and (CDN_nD_nE_nSI, CDN, nD, nE, nSI);
    and (CDN_D_E_SE, CDN, D, E, SE);
    and (CDN_nD_E_SE, CDN, nD, E, SE);
    and (CDN_D_nE_SE, CDN, D, nE, SE);
    and (CDN_nD_nE_SE, CDN, nD, nE, SE);
    and (D_E_SE_SI, D, E, SE, SI);
    and (D_E_nSE_SI, D, E, nSE, SI);
    and (D_E_nSE_nSI, D, E, nSE, nSI);
    and (nD_E_SE_SI, nD, E, SE, SI);
    and (D_nE_SE_SI, D, nE, SE, SI);
    and (nD_nE_SE_SI, nD, nE, SE, SI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
    and  (D_check, CDN_i, E_d, SE_int_not);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
    and  (D_check, CDN_i, E, SE_int_not);
  `endif
  and  (E_check, CDN_i, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (negedge CDN &&& CP_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_E_SE_SI_SDFCHK, posedge CP &&& D_E_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_E_nSE_SI_SDFCHK, posedge CP &&& D_E_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_E_nSE_nSI_SDFCHK, posedge CP &&& D_E_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_E_SE_SI_SDFCHK, posedge CP &&& nD_E_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nE_SE_SI_SDFCHK, posedge CP &&& D_nE_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_nE_SE_SI_SDFCHK, posedge CP &&& nD_nE_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_E_SE_SI_SDFCHK, posedge CP &&& D_E_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_E_nSE_SI_SDFCHK, posedge CP &&& D_E_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_E_nSE_nSI_SDFCHK, posedge CP &&& D_E_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_E_SE_SI_SDFCHK, posedge CP &&& nD_E_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nE_SE_SI_SDFCHK, posedge CP &&& D_nE_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_nE_SE_SI_SDFCHK, posedge CP &&& nD_nE_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_E_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_E_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_E_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_E_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nE_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_nE_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_E_SE_SI_SDFCHK, posedge CP &&& D_E_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_E_nSE_SI_SDFCHK, posedge CP &&& D_E_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_E_nSE_nSI_SDFCHK, posedge CP &&& D_E_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_E_SE_SI_SDFCHK, posedge CP &&& nD_E_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nE_SE_SI_SDFCHK, posedge CP &&& D_nE_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_nE_SE_SI_SDFCHK, posedge CP &&& nD_nE_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_E_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_E_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_E_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_E_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nE_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_nE_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFCNQD2 (E, SE, CP, SI, D, CDN, Q);
    input E, SE, CP, SI, D, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire E_d, SE_d, CP_d, SI_d, D_d;
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_E_SE_SI_SDFCHK, CP_D_E_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_E_SE_nSI_SDFCHK, CP_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_E_nSE_SI_SDFCHK, CP_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_E_nSE_nSI_SDFCHK, CP_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_E_SE_SI_SDFCHK, CP_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_E_SE_nSI_SDFCHK, CP_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_E_nSE_SI_SDFCHK, CP_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_E_nSE_nSI_SDFCHK, CP_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nE_SE_SI_SDFCHK, CP_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_nE_SE_nSI_SDFCHK, CP_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nE_nSE_SI_SDFCHK, CP_D_nE_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nE_nSE_nSI_SDFCHK, CP_D_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nE_SE_SI_SDFCHK, CP_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nE_SE_nSI_SDFCHK, CP_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nE_nSE_SI_SDFCHK, CP_nD_nE_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nE_nSE_nSI_SDFCHK, CP_nD_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_E_SE_SI_SDFCHK, nCP_D_E_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_E_SE_nSI_SDFCHK, nCP_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_E_nSE_SI_SDFCHK, nCP_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_E_nSE_nSI_SDFCHK, nCP_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_E_SE_SI_SDFCHK, nCP_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_E_SE_nSI_SDFCHK, nCP_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_E_nSE_SI_SDFCHK, nCP_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_E_nSE_nSI_SDFCHK, nCP_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nE_SE_SI_SDFCHK, nCP_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nE_SE_nSI_SDFCHK, nCP_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nE_nSE_SI_SDFCHK, nCP_D_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nE_nSE_nSI_SDFCHK, nCP_D_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nE_SE_SI_SDFCHK, nCP_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nE_SE_nSI_SDFCHK, nCP_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nE_nSE_SI_SDFCHK, nCP_nD_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nE_nSE_nSI_SDFCHK, nCP_nD_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_E_SE_SI_SDFCHK, CDN_D_E_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_E_nSE_SI_SDFCHK, CDN_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_E_nSE_nSI_SDFCHK, CDN_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_E_SE_SI_SDFCHK, CDN_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nE_SE_SI_SDFCHK, CDN_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SE_SI_SDFCHK, CDN_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_E_SE_nSI_SDFCHK, CDN_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_E_SE_nSI_SDFCHK, CDN_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_E_nSE_SI_SDFCHK, CDN_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_E_nSE_nSI_SDFCHK, CDN_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_nE_SE_nSI_SDFCHK, CDN_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SE_nSI_SDFCHK, CDN_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_E_nSE_SI_SDFCHK, CDN_E_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_E_nSE_nSI_SDFCHK, CDN_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_nE_SI_SDFCHK, CDN_D_nE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SI_SDFCHK, CDN_nD_nE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_E_SI_SDFCHK, CDN_nD_E_SI, 1'b1);
    tsmc_xbuf (CDN_D_E_nSI_SDFCHK, CDN_D_E_nSI, 1'b1);
    tsmc_xbuf (CDN_D_nE_nSI_SDFCHK, CDN_D_nE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nE_nSI_SDFCHK, CDN_nD_nE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_E_SE_SDFCHK, CDN_D_E_SE, 1'b1);
    tsmc_xbuf (CDN_nD_E_SE_SDFCHK, CDN_nD_E_SE, 1'b1);
    tsmc_xbuf (CDN_D_nE_SE_SDFCHK, CDN_D_nE_SE, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SE_SDFCHK, CDN_nD_nE_SE, 1'b1);
    tsmc_xbuf (D_E_SE_SI_SDFCHK, D_E_SE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_SI_SDFCHK, D_E_nSE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_nSI_SDFCHK, D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_E_SE_SI_SDFCHK, nD_E_SE_SI, 1'b1);
    tsmc_xbuf (D_nE_SE_SI_SDFCHK, D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SE_SI_SDFCHK, nD_nE_SE_SI, 1'b1);
  `endif

    not (nE, E);
    not (nSE, SE);
    not (nCP, CP);
    not (nSI, SI);
    not (nD, D);
    and (CP_D_E_SE_SI, CP, D, E, SE, SI);
    and (CP_D_E_SE_nSI, CP, D, E, SE, nSI);
    and (CP_D_E_nSE_SI, CP, D, E, nSE, SI);
    and (CP_D_E_nSE_nSI, CP, D, E, nSE, nSI);
    and (CP_nD_E_SE_SI, CP, nD, E, SE, SI);
    and (CP_nD_E_SE_nSI, CP, nD, E, SE, nSI);
    and (CP_nD_E_nSE_SI, CP, nD, E, nSE, SI);
    and (CP_nD_E_nSE_nSI, CP, nD, E, nSE, nSI);
    and (CP_D_nE_SE_SI, CP, D, nE, SE, SI);
    and (CP_D_nE_SE_nSI, CP, D, nE, SE, nSI);
    and (CP_D_nE_nSE_SI, CP, D, nE, nSE, SI);
    and (CP_D_nE_nSE_nSI, CP, D, nE, nSE, nSI);
    and (CP_nD_nE_SE_SI, CP, nD, nE, SE, SI);
    and (CP_nD_nE_SE_nSI, CP, nD, nE, SE, nSI);
    and (CP_nD_nE_nSE_SI, CP, nD, nE, nSE, SI);
    and (CP_nD_nE_nSE_nSI, CP, nD, nE, nSE, nSI);
    and (nCP_D_E_SE_SI, nCP, D, E, SE, SI);
    and (nCP_D_E_SE_nSI, nCP, D, E, SE, nSI);
    and (nCP_D_E_nSE_SI, nCP, D, E, nSE, SI);
    and (nCP_D_E_nSE_nSI, nCP, D, E, nSE, nSI);
    and (nCP_nD_E_SE_SI, nCP, nD, E, SE, SI);
    and (nCP_nD_E_SE_nSI, nCP, nD, E, SE, nSI);
    and (nCP_nD_E_nSE_SI, nCP, nD, E, nSE, SI);
    and (nCP_nD_E_nSE_nSI, nCP, nD, E, nSE, nSI);
    and (nCP_D_nE_SE_SI, nCP, D, nE, SE, SI);
    and (nCP_D_nE_SE_nSI, nCP, D, nE, SE, nSI);
    and (nCP_D_nE_nSE_SI, nCP, D, nE, nSE, SI);
    and (nCP_D_nE_nSE_nSI, nCP, D, nE, nSE, nSI);
    and (nCP_nD_nE_SE_SI, nCP, nD, nE, SE, SI);
    and (nCP_nD_nE_SE_nSI, nCP, nD, nE, SE, nSI);
    and (nCP_nD_nE_nSE_SI, nCP, nD, nE, nSE, SI);
    and (nCP_nD_nE_nSE_nSI, nCP, nD, nE, nSE, nSI);
    and (CDN_D_E_SE_SI, CDN, D, E, SE, SI);
    and (CDN_D_E_nSE_SI, CDN, D, E, nSE, SI);
    and (CDN_D_E_nSE_nSI, CDN, D, E, nSE, nSI);
    and (CDN_nD_E_SE_SI, CDN, nD, E, SE, SI);
    and (CDN_D_nE_SE_SI, CDN, D, nE, SE, SI);
    and (CDN_nD_nE_SE_SI, CDN, nD, nE, SE, SI);
    and (CDN_D_E_SE_nSI, CDN, D, E, SE, nSI);
    and (CDN_nD_E_SE_nSI, CDN, nD, E, SE, nSI);
    and (CDN_nD_E_nSE_SI, CDN, nD, E, nSE, SI);
    and (CDN_nD_E_nSE_nSI, CDN, nD, E, nSE, nSI);
    and (CDN_D_nE_SE_nSI, CDN, D, nE, SE, nSI);
    and (CDN_nD_nE_SE_nSI, CDN, nD, nE, SE, nSI);
    and (CDN_E_nSE_SI, CDN, E, nSE, SI);
    and (CDN_E_nSE_nSI, CDN, E, nSE, nSI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_D_nE_SI, CDN, D, nE, SI);
    and (CDN_nD_nE_SI, CDN, nD, nE, SI);
    and (CDN_nD_E_SI, CDN, nD, E, SI);
    and (CDN_D_E_nSI, CDN, D, E, nSI);
    and (CDN_D_nE_nSI, CDN, D, nE, nSI);
    and (CDN_nD_nE_nSI, CDN, nD, nE, nSI);
    and (CDN_D_E_SE, CDN, D, E, SE);
    and (CDN_nD_E_SE, CDN, nD, E, SE);
    and (CDN_D_nE_SE, CDN, D, nE, SE);
    and (CDN_nD_nE_SE, CDN, nD, nE, SE);
    and (D_E_SE_SI, D, E, SE, SI);
    and (D_E_nSE_SI, D, E, nSE, SI);
    and (D_E_nSE_nSI, D, E, nSE, nSI);
    and (nD_E_SE_SI, nD, E, SE, SI);
    and (D_nE_SE_SI, D, nE, SE, SI);
    and (nD_nE_SE_SI, nD, nE, SE, SI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
    and  (D_check, CDN_i, E_d, SE_int_not);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
    and  (D_check, CDN_i, E, SE_int_not);
  `endif
  and  (E_check, CDN_i, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (negedge CDN &&& CP_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_E_SE_SI_SDFCHK, posedge CP &&& D_E_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_E_nSE_SI_SDFCHK, posedge CP &&& D_E_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_E_nSE_nSI_SDFCHK, posedge CP &&& D_E_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_E_SE_SI_SDFCHK, posedge CP &&& nD_E_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nE_SE_SI_SDFCHK, posedge CP &&& D_nE_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_nE_SE_SI_SDFCHK, posedge CP &&& nD_nE_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_E_SE_SI_SDFCHK, posedge CP &&& D_E_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_E_nSE_SI_SDFCHK, posedge CP &&& D_E_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_E_nSE_nSI_SDFCHK, posedge CP &&& D_E_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_E_SE_SI_SDFCHK, posedge CP &&& nD_E_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nE_SE_SI_SDFCHK, posedge CP &&& D_nE_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_nE_SE_SI_SDFCHK, posedge CP &&& nD_nE_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_E_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_E_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_E_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_E_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nE_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_nE_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_E_SE_SI_SDFCHK, posedge CP &&& D_E_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_E_nSE_SI_SDFCHK, posedge CP &&& D_E_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_E_nSE_nSI_SDFCHK, posedge CP &&& D_E_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_E_SE_SI_SDFCHK, posedge CP &&& nD_E_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nE_SE_SI_SDFCHK, posedge CP &&& D_nE_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_nE_SE_SI_SDFCHK, posedge CP &&& nD_nE_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_E_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_E_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_E_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_E_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nE_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_nE_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFCNQD4 (E, SE, CP, SI, D, CDN, Q);
    input E, SE, CP, SI, D, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire E_d, SE_d, CP_d, SI_d, D_d;
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_E_SE_SI_SDFCHK, CP_D_E_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_E_SE_nSI_SDFCHK, CP_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_E_nSE_SI_SDFCHK, CP_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_E_nSE_nSI_SDFCHK, CP_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_E_SE_SI_SDFCHK, CP_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_E_SE_nSI_SDFCHK, CP_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_E_nSE_SI_SDFCHK, CP_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_E_nSE_nSI_SDFCHK, CP_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nE_SE_SI_SDFCHK, CP_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_nE_SE_nSI_SDFCHK, CP_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nE_nSE_SI_SDFCHK, CP_D_nE_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nE_nSE_nSI_SDFCHK, CP_D_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nE_SE_SI_SDFCHK, CP_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nE_SE_nSI_SDFCHK, CP_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nE_nSE_SI_SDFCHK, CP_nD_nE_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nE_nSE_nSI_SDFCHK, CP_nD_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_E_SE_SI_SDFCHK, nCP_D_E_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_E_SE_nSI_SDFCHK, nCP_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_E_nSE_SI_SDFCHK, nCP_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_E_nSE_nSI_SDFCHK, nCP_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_E_SE_SI_SDFCHK, nCP_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_E_SE_nSI_SDFCHK, nCP_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_E_nSE_SI_SDFCHK, nCP_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_E_nSE_nSI_SDFCHK, nCP_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nE_SE_SI_SDFCHK, nCP_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nE_SE_nSI_SDFCHK, nCP_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nE_nSE_SI_SDFCHK, nCP_D_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nE_nSE_nSI_SDFCHK, nCP_D_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nE_SE_SI_SDFCHK, nCP_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nE_SE_nSI_SDFCHK, nCP_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nE_nSE_SI_SDFCHK, nCP_nD_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nE_nSE_nSI_SDFCHK, nCP_nD_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_E_SE_SI_SDFCHK, CDN_D_E_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_E_nSE_SI_SDFCHK, CDN_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_E_nSE_nSI_SDFCHK, CDN_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_E_SE_SI_SDFCHK, CDN_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nE_SE_SI_SDFCHK, CDN_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SE_SI_SDFCHK, CDN_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_E_SE_nSI_SDFCHK, CDN_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_E_SE_nSI_SDFCHK, CDN_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_E_nSE_SI_SDFCHK, CDN_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_E_nSE_nSI_SDFCHK, CDN_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_nE_SE_nSI_SDFCHK, CDN_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SE_nSI_SDFCHK, CDN_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_E_nSE_SI_SDFCHK, CDN_E_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_E_nSE_nSI_SDFCHK, CDN_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_nE_SI_SDFCHK, CDN_D_nE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SI_SDFCHK, CDN_nD_nE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_E_SI_SDFCHK, CDN_nD_E_SI, 1'b1);
    tsmc_xbuf (CDN_D_E_nSI_SDFCHK, CDN_D_E_nSI, 1'b1);
    tsmc_xbuf (CDN_D_nE_nSI_SDFCHK, CDN_D_nE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nE_nSI_SDFCHK, CDN_nD_nE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_E_SE_SDFCHK, CDN_D_E_SE, 1'b1);
    tsmc_xbuf (CDN_nD_E_SE_SDFCHK, CDN_nD_E_SE, 1'b1);
    tsmc_xbuf (CDN_D_nE_SE_SDFCHK, CDN_D_nE_SE, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SE_SDFCHK, CDN_nD_nE_SE, 1'b1);
    tsmc_xbuf (D_E_SE_SI_SDFCHK, D_E_SE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_SI_SDFCHK, D_E_nSE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_nSI_SDFCHK, D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_E_SE_SI_SDFCHK, nD_E_SE_SI, 1'b1);
    tsmc_xbuf (D_nE_SE_SI_SDFCHK, D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SE_SI_SDFCHK, nD_nE_SE_SI, 1'b1);
  `endif

    not (nE, E);
    not (nSE, SE);
    not (nCP, CP);
    not (nSI, SI);
    not (nD, D);
    and (CP_D_E_SE_SI, CP, D, E, SE, SI);
    and (CP_D_E_SE_nSI, CP, D, E, SE, nSI);
    and (CP_D_E_nSE_SI, CP, D, E, nSE, SI);
    and (CP_D_E_nSE_nSI, CP, D, E, nSE, nSI);
    and (CP_nD_E_SE_SI, CP, nD, E, SE, SI);
    and (CP_nD_E_SE_nSI, CP, nD, E, SE, nSI);
    and (CP_nD_E_nSE_SI, CP, nD, E, nSE, SI);
    and (CP_nD_E_nSE_nSI, CP, nD, E, nSE, nSI);
    and (CP_D_nE_SE_SI, CP, D, nE, SE, SI);
    and (CP_D_nE_SE_nSI, CP, D, nE, SE, nSI);
    and (CP_D_nE_nSE_SI, CP, D, nE, nSE, SI);
    and (CP_D_nE_nSE_nSI, CP, D, nE, nSE, nSI);
    and (CP_nD_nE_SE_SI, CP, nD, nE, SE, SI);
    and (CP_nD_nE_SE_nSI, CP, nD, nE, SE, nSI);
    and (CP_nD_nE_nSE_SI, CP, nD, nE, nSE, SI);
    and (CP_nD_nE_nSE_nSI, CP, nD, nE, nSE, nSI);
    and (nCP_D_E_SE_SI, nCP, D, E, SE, SI);
    and (nCP_D_E_SE_nSI, nCP, D, E, SE, nSI);
    and (nCP_D_E_nSE_SI, nCP, D, E, nSE, SI);
    and (nCP_D_E_nSE_nSI, nCP, D, E, nSE, nSI);
    and (nCP_nD_E_SE_SI, nCP, nD, E, SE, SI);
    and (nCP_nD_E_SE_nSI, nCP, nD, E, SE, nSI);
    and (nCP_nD_E_nSE_SI, nCP, nD, E, nSE, SI);
    and (nCP_nD_E_nSE_nSI, nCP, nD, E, nSE, nSI);
    and (nCP_D_nE_SE_SI, nCP, D, nE, SE, SI);
    and (nCP_D_nE_SE_nSI, nCP, D, nE, SE, nSI);
    and (nCP_D_nE_nSE_SI, nCP, D, nE, nSE, SI);
    and (nCP_D_nE_nSE_nSI, nCP, D, nE, nSE, nSI);
    and (nCP_nD_nE_SE_SI, nCP, nD, nE, SE, SI);
    and (nCP_nD_nE_SE_nSI, nCP, nD, nE, SE, nSI);
    and (nCP_nD_nE_nSE_SI, nCP, nD, nE, nSE, SI);
    and (nCP_nD_nE_nSE_nSI, nCP, nD, nE, nSE, nSI);
    and (CDN_D_E_SE_SI, CDN, D, E, SE, SI);
    and (CDN_D_E_nSE_SI, CDN, D, E, nSE, SI);
    and (CDN_D_E_nSE_nSI, CDN, D, E, nSE, nSI);
    and (CDN_nD_E_SE_SI, CDN, nD, E, SE, SI);
    and (CDN_D_nE_SE_SI, CDN, D, nE, SE, SI);
    and (CDN_nD_nE_SE_SI, CDN, nD, nE, SE, SI);
    and (CDN_D_E_SE_nSI, CDN, D, E, SE, nSI);
    and (CDN_nD_E_SE_nSI, CDN, nD, E, SE, nSI);
    and (CDN_nD_E_nSE_SI, CDN, nD, E, nSE, SI);
    and (CDN_nD_E_nSE_nSI, CDN, nD, E, nSE, nSI);
    and (CDN_D_nE_SE_nSI, CDN, D, nE, SE, nSI);
    and (CDN_nD_nE_SE_nSI, CDN, nD, nE, SE, nSI);
    and (CDN_E_nSE_SI, CDN, E, nSE, SI);
    and (CDN_E_nSE_nSI, CDN, E, nSE, nSI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_D_nE_SI, CDN, D, nE, SI);
    and (CDN_nD_nE_SI, CDN, nD, nE, SI);
    and (CDN_nD_E_SI, CDN, nD, E, SI);
    and (CDN_D_E_nSI, CDN, D, E, nSI);
    and (CDN_D_nE_nSI, CDN, D, nE, nSI);
    and (CDN_nD_nE_nSI, CDN, nD, nE, nSI);
    and (CDN_D_E_SE, CDN, D, E, SE);
    and (CDN_nD_E_SE, CDN, nD, E, SE);
    and (CDN_D_nE_SE, CDN, D, nE, SE);
    and (CDN_nD_nE_SE, CDN, nD, nE, SE);
    and (D_E_SE_SI, D, E, SE, SI);
    and (D_E_nSE_SI, D, E, nSE, SI);
    and (D_E_nSE_nSI, D, E, nSE, nSI);
    and (nD_E_SE_SI, nD, E, SE, SI);
    and (D_nE_SE_SI, D, nE, SE, SI);
    and (nD_nE_SE_SI, nD, nE, SE, SI);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
    and  (D_check, CDN_i, E_d, SE_int_not);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
    and  (D_check, CDN_i, E, SE_int_not);
  `endif
  and  (E_check, CDN_i, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && E == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (negedge CDN &&& CP_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_E_SE_SI_SDFCHK, posedge CP &&& D_E_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_E_nSE_SI_SDFCHK, posedge CP &&& D_E_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_E_nSE_nSI_SDFCHK, posedge CP &&& D_E_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_E_SE_SI_SDFCHK, posedge CP &&& nD_E_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nE_SE_SI_SDFCHK, posedge CP &&& D_nE_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_nE_SE_SI_SDFCHK, posedge CP &&& nD_nE_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_E_SE_SI_SDFCHK, posedge CP &&& D_E_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_E_nSE_SI_SDFCHK, posedge CP &&& D_E_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_E_nSE_nSI_SDFCHK, posedge CP &&& D_E_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_E_SE_SI_SDFCHK, posedge CP &&& nD_E_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nE_SE_SI_SDFCHK, posedge CP &&& D_nE_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_nE_SE_SI_SDFCHK, posedge CP &&& nD_nE_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_E_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_E_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_E_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_E_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nE_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_nE_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_E_SE_SI_SDFCHK, posedge CP &&& D_E_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_E_nSE_SI_SDFCHK, posedge CP &&& D_E_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_E_nSE_nSI_SDFCHK, posedge CP &&& D_E_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_E_SE_SI_SDFCHK, posedge CP &&& nD_E_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nE_SE_SI_SDFCHK, posedge CP &&& D_nE_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_nE_SE_SI_SDFCHK, posedge CP &&& nD_nE_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_E_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_E_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_E_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_E_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nE_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_nE_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFD0 (E, SE, CP, SI, D, Q, QN);
    input E, SE, CP, SI, D;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire E_d, SE_d, CP_d, SI_d, D_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_E_SE_SI_SDFCHK, D_E_SE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_SI_SDFCHK, D_E_nSE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_nSI_SDFCHK, D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_E_SE_SI_SDFCHK, nD_E_SE_SI, 1'b1);
    tsmc_xbuf (D_nE_SE_SI_SDFCHK, D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SE_SI_SDFCHK, nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (D_E_SE_nSI_SDFCHK, D_E_SE_nSI, 1'b1);
    tsmc_xbuf (nD_E_SE_nSI_SDFCHK, nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (nD_E_nSE_SI_SDFCHK, nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (nD_E_nSE_nSI_SDFCHK, nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nE_SE_nSI_SDFCHK, D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_SE_nSI_SDFCHK, nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (E_nSE_SI_SDFCHK, E_nSE_SI, 1'b1);
    tsmc_xbuf (E_nSE_nSI_SDFCHK, E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nE_SI_SDFCHK, D_nE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SI_SDFCHK, nD_nE_SI, 1'b1);
    tsmc_xbuf (nD_E_SI_SDFCHK, nD_E_SI, 1'b1);
    tsmc_xbuf (D_E_nSI_SDFCHK, D_E_nSI, 1'b1);
    tsmc_xbuf (D_nE_nSI_SDFCHK, D_nE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_nSI_SDFCHK, nD_nE_nSI, 1'b1);
    tsmc_xbuf (D_E_SE_SDFCHK, D_E_SE, 1'b1);
    tsmc_xbuf (D_nE_SE_SDFCHK, D_nE_SE, 1'b1);
    tsmc_xbuf (nD_nE_SE_SDFCHK, nD_nE_SE, 1'b1);
    tsmc_xbuf (nD_E_SE_SDFCHK, nD_E_SE, 1'b1);
  `endif

    not (nE, E);
    not (nSE, SE);
    not (nSI, SI);
    not (nD, D);
    and (D_E_SE_SI, D, E, SE, SI);
    and (D_E_nSE_SI, D, E, nSE, SI);
    and (D_E_nSE_nSI, D, E, nSE, nSI);
    and (nD_E_SE_SI, nD, E, SE, SI);
    and (D_nE_SE_SI, D, nE, SE, SI);
    and (nD_nE_SE_SI, nD, nE, SE, SI);
    and (D_E_SE_nSI, D, E, SE, nSI);
    and (nD_E_SE_nSI, nD, E, SE, nSI);
    and (nD_E_nSE_SI, nD, E, nSE, SI);
    and (nD_E_nSE_nSI, nD, E, nSE, nSI);
    and (D_nE_SE_nSI, D, nE, SE, nSI);
    and (nD_nE_SE_nSI, nD, nE, SE, nSI);
    and (E_nSE_SI, E, nSE, SI);
    and (E_nSE_nSI, E, nSE, nSI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (D_nE_SI, D, nE, SI);
    and (nD_nE_SI, nD, nE, SI);
    and (nD_E_SI, nD, E, SI);
    and (D_E_nSI, D, E, nSI);
    and (D_nE_nSI, D, nE, nSI);
    and (nD_nE_nSI, nD, nE, nSI);
    and (D_E_SE, D, E, SE);
    and (D_nE_SE, D, nE, SE);
    and (nD_nE_SE, nD, nE, SE);
    and (nD_E_SE, nD, E, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFD1 (E, SE, CP, SI, D, Q, QN);
    input E, SE, CP, SI, D;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire E_d, SE_d, CP_d, SI_d, D_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_E_SE_SI_SDFCHK, D_E_SE_SI, 1'b1);
    tsmc_xbuf (D_nE_SE_SI_SDFCHK, D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nD_E_SE_SI_SDFCHK, nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SE_SI_SDFCHK, nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_SI_SDFCHK, D_E_nSE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_nSI_SDFCHK, D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_E_SE_nSI_SDFCHK, D_E_SE_nSI, 1'b1);
    tsmc_xbuf (D_nE_SE_nSI_SDFCHK, D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nD_E_SE_nSI_SDFCHK, nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_SE_nSI_SDFCHK, nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nD_E_nSE_SI_SDFCHK, nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (nD_E_nSE_nSI_SDFCHK, nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (E_nSE_SI_SDFCHK, E_nSE_SI, 1'b1);
    tsmc_xbuf (E_nSE_nSI_SDFCHK, E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nE_SI_SDFCHK, D_nE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SI_SDFCHK, nD_nE_SI, 1'b1);
    tsmc_xbuf (nD_E_SI_SDFCHK, nD_E_SI, 1'b1);
    tsmc_xbuf (D_E_nSI_SDFCHK, D_E_nSI, 1'b1);
    tsmc_xbuf (D_nE_nSI_SDFCHK, D_nE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_nSI_SDFCHK, nD_nE_nSI, 1'b1);
    tsmc_xbuf (D_E_SE_SDFCHK, D_E_SE, 1'b1);
    tsmc_xbuf (nD_E_SE_SDFCHK, nD_E_SE, 1'b1);
    tsmc_xbuf (D_nE_SE_SDFCHK, D_nE_SE, 1'b1);
    tsmc_xbuf (nD_nE_SE_SDFCHK, nD_nE_SE, 1'b1);
  `endif

    not (nE, E);
    not (nSE, SE);
    not (nSI, SI);
    not (nD, D);
    and (D_E_SE_SI, D, E, SE, SI);
    and (D_nE_SE_SI, D, nE, SE, SI);
    and (nD_E_SE_SI, nD, E, SE, SI);
    and (nD_nE_SE_SI, nD, nE, SE, SI);
    and (D_E_nSE_SI, D, E, nSE, SI);
    and (D_E_nSE_nSI, D, E, nSE, nSI);
    and (D_E_SE_nSI, D, E, SE, nSI);
    and (D_nE_SE_nSI, D, nE, SE, nSI);
    and (nD_E_SE_nSI, nD, E, SE, nSI);
    and (nD_nE_SE_nSI, nD, nE, SE, nSI);
    and (nD_E_nSE_SI, nD, E, nSE, SI);
    and (nD_E_nSE_nSI, nD, E, nSE, nSI);
    and (E_nSE_SI, E, nSE, SI);
    and (E_nSE_nSI, E, nSE, nSI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (D_nE_SI, D, nE, SI);
    and (nD_nE_SI, nD, nE, SI);
    and (nD_E_SI, nD, E, SI);
    and (D_E_nSI, D, E, nSI);
    and (D_nE_nSI, D, nE, nSI);
    and (nD_nE_nSI, nD, nE, nSI);
    and (D_E_SE, D, E, SE);
    and (nD_E_SE, nD, E, SE);
    and (D_nE_SE, D, nE, SE);
    and (nD_nE_SE, nD, nE, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFD2 (E, SE, CP, SI, D, Q, QN);
    input E, SE, CP, SI, D;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire E_d, SE_d, CP_d, SI_d, D_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_E_SE_SI_SDFCHK, D_E_SE_SI, 1'b1);
    tsmc_xbuf (D_nE_SE_SI_SDFCHK, D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nD_E_SE_SI_SDFCHK, nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SE_SI_SDFCHK, nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_SI_SDFCHK, D_E_nSE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_nSI_SDFCHK, D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_E_SE_nSI_SDFCHK, D_E_SE_nSI, 1'b1);
    tsmc_xbuf (D_nE_SE_nSI_SDFCHK, D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nD_E_SE_nSI_SDFCHK, nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_SE_nSI_SDFCHK, nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nD_E_nSE_SI_SDFCHK, nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (nD_E_nSE_nSI_SDFCHK, nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (E_nSE_SI_SDFCHK, E_nSE_SI, 1'b1);
    tsmc_xbuf (E_nSE_nSI_SDFCHK, E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nE_SI_SDFCHK, D_nE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SI_SDFCHK, nD_nE_SI, 1'b1);
    tsmc_xbuf (nD_E_SI_SDFCHK, nD_E_SI, 1'b1);
    tsmc_xbuf (D_E_nSI_SDFCHK, D_E_nSI, 1'b1);
    tsmc_xbuf (D_nE_nSI_SDFCHK, D_nE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_nSI_SDFCHK, nD_nE_nSI, 1'b1);
    tsmc_xbuf (D_E_SE_SDFCHK, D_E_SE, 1'b1);
    tsmc_xbuf (nD_E_SE_SDFCHK, nD_E_SE, 1'b1);
    tsmc_xbuf (D_nE_SE_SDFCHK, D_nE_SE, 1'b1);
    tsmc_xbuf (nD_nE_SE_SDFCHK, nD_nE_SE, 1'b1);
  `endif

    not (nE, E);
    not (nSE, SE);
    not (nSI, SI);
    not (nD, D);
    and (D_E_SE_SI, D, E, SE, SI);
    and (D_nE_SE_SI, D, nE, SE, SI);
    and (nD_E_SE_SI, nD, E, SE, SI);
    and (nD_nE_SE_SI, nD, nE, SE, SI);
    and (D_E_nSE_SI, D, E, nSE, SI);
    and (D_E_nSE_nSI, D, E, nSE, nSI);
    and (D_E_SE_nSI, D, E, SE, nSI);
    and (D_nE_SE_nSI, D, nE, SE, nSI);
    and (nD_E_SE_nSI, nD, E, SE, nSI);
    and (nD_nE_SE_nSI, nD, nE, SE, nSI);
    and (nD_E_nSE_SI, nD, E, nSE, SI);
    and (nD_E_nSE_nSI, nD, E, nSE, nSI);
    and (E_nSE_SI, E, nSE, SI);
    and (E_nSE_nSI, E, nSE, nSI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (D_nE_SI, D, nE, SI);
    and (nD_nE_SI, nD, nE, SI);
    and (nD_E_SI, nD, E, SI);
    and (D_E_nSI, D, E, nSI);
    and (D_nE_nSI, D, nE, nSI);
    and (nD_nE_nSI, nD, nE, nSI);
    and (D_E_SE, D, E, SE);
    and (nD_E_SE, nD, E, SE);
    and (D_nE_SE, D, nE, SE);
    and (nD_nE_SE, nD, nE, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFD4 (E, SE, CP, SI, D, Q, QN);
    input E, SE, CP, SI, D;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire E_d, SE_d, CP_d, SI_d, D_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_E_SE_SI_SDFCHK, D_E_SE_SI, 1'b1);
    tsmc_xbuf (D_nE_SE_SI_SDFCHK, D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nD_E_SE_SI_SDFCHK, nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SE_SI_SDFCHK, nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_SI_SDFCHK, D_E_nSE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_nSI_SDFCHK, D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_E_SE_nSI_SDFCHK, D_E_SE_nSI, 1'b1);
    tsmc_xbuf (D_nE_SE_nSI_SDFCHK, D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nD_E_SE_nSI_SDFCHK, nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_SE_nSI_SDFCHK, nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nD_E_nSE_SI_SDFCHK, nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (nD_E_nSE_nSI_SDFCHK, nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (E_nSE_SI_SDFCHK, E_nSE_SI, 1'b1);
    tsmc_xbuf (E_nSE_nSI_SDFCHK, E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nE_SI_SDFCHK, D_nE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SI_SDFCHK, nD_nE_SI, 1'b1);
    tsmc_xbuf (nD_E_SI_SDFCHK, nD_E_SI, 1'b1);
    tsmc_xbuf (D_E_nSI_SDFCHK, D_E_nSI, 1'b1);
    tsmc_xbuf (D_nE_nSI_SDFCHK, D_nE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_nSI_SDFCHK, nD_nE_nSI, 1'b1);
    tsmc_xbuf (D_E_SE_SDFCHK, D_E_SE, 1'b1);
    tsmc_xbuf (nD_E_SE_SDFCHK, nD_E_SE, 1'b1);
    tsmc_xbuf (D_nE_SE_SDFCHK, D_nE_SE, 1'b1);
    tsmc_xbuf (nD_nE_SE_SDFCHK, nD_nE_SE, 1'b1);
  `endif

    not (nE, E);
    not (nSE, SE);
    not (nSI, SI);
    not (nD, D);
    and (D_E_SE_SI, D, E, SE, SI);
    and (D_nE_SE_SI, D, nE, SE, SI);
    and (nD_E_SE_SI, nD, E, SE, SI);
    and (nD_nE_SE_SI, nD, nE, SE, SI);
    and (D_E_nSE_SI, D, E, nSE, SI);
    and (D_E_nSE_nSI, D, E, nSE, nSI);
    and (D_E_SE_nSI, D, E, SE, nSI);
    and (D_nE_SE_nSI, D, nE, SE, nSI);
    and (nD_E_SE_nSI, nD, E, SE, nSI);
    and (nD_nE_SE_nSI, nD, nE, SE, nSI);
    and (nD_E_nSE_SI, nD, E, nSE, SI);
    and (nD_E_nSE_nSI, nD, E, nSE, nSI);
    and (E_nSE_SI, E, nSE, SI);
    and (E_nSE_nSI, E, nSE, nSI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (D_nE_SI, D, nE, SI);
    and (nD_nE_SI, nD, nE, SI);
    and (nD_E_SI, nD, E, SI);
    and (D_E_nSI, D, E, nSI);
    and (D_nE_nSI, D, nE, nSI);
    and (nD_nE_nSI, nD, nE, nSI);
    and (D_E_SE, D, E, SE);
    and (nD_E_SE, nD, E, SE);
    and (D_nE_SE, D, nE, SE);
    and (nD_nE_SE, nD, nE, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFKCND0 (SI, D, E, SE, CP, CN, Q, QN);
    input SI, D, SE, CP, CN, E;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d, E_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        and (D2, CN_d, D1);
        tsmc_mux (D3, D2, SI_d, SE_d);
        tsmc_dff (Q_buf, D3, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        and (D2, CN, D1);
        tsmc_mux (D3, D2, SI, SE);
        tsmc_dff (Q_buf, D3, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_E_SE_SI_SDFCHK, CN_D_E_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_E_nSE_SI_SDFCHK, CN_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (CN_D_E_nSE_nSI_SDFCHK, CN_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_E_SE_SI_SDFCHK, CN_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nCN_D_E_SE_SI_SDFCHK, nCN_D_E_SE_SI, 1'b1);
    tsmc_xbuf (nCN_D_nE_SE_SI_SDFCHK, nCN_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_E_SE_SI_SDFCHK, nCN_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SE_SI_SDFCHK, nCN_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_nE_SE_SI_SDFCHK, CN_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nE_SE_SI_SDFCHK, CN_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_E_SE_nSI_SDFCHK, CN_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_E_SE_nSI_SDFCHK, CN_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_E_nSE_SI_SDFCHK, CN_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_E_nSE_nSI_SDFCHK, CN_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_E_SE_nSI_SDFCHK, nCN_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_E_nSE_SI_SDFCHK, nCN_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_D_E_nSE_nSI_SDFCHK, nCN_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_nE_SE_nSI_SDFCHK, nCN_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_nE_nSE_SI_SDFCHK, nCN_D_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_D_nE_nSE_nSI_SDFCHK, nCN_D_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_E_SE_nSI_SDFCHK, nCN_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_E_nSE_SI_SDFCHK, nCN_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_E_nSE_nSI_SDFCHK, nCN_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SE_nSI_SDFCHK, nCN_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_nSE_SI_SDFCHK, nCN_nD_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_nSE_nSI_SDFCHK, nCN_nD_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_D_nE_SE_nSI_SDFCHK, CN_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nE_SE_nSI_SDFCHK, CN_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (D_E_nSE_SI_SDFCHK, D_E_nSE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_nSI_SDFCHK, D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nE_nSE_SI_SDFCHK, D_nE_nSE_SI, 1'b1);
    tsmc_xbuf (D_nE_nSE_nSI_SDFCHK, D_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_nSE_SI_SDFCHK, nD_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nE_nSE_nSI_SDFCHK, nD_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_E_nSE_SI_SDFCHK, CN_E_nSE_SI, 1'b1);
    tsmc_xbuf (CN_E_nSE_nSI_SDFCHK, CN_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SDFCHK, CN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SDFCHK, CN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_D_nE_SI_SDFCHK, CN_D_nE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nE_SI_SDFCHK, CN_nD_nE_SI, 1'b1);
    tsmc_xbuf (CN_nD_E_SI_SDFCHK, CN_nD_E_SI, 1'b1);
    tsmc_xbuf (nCN_D_E_SI_SDFCHK, nCN_D_E_SI, 1'b1);
    tsmc_xbuf (nCN_D_nE_SI_SDFCHK, nCN_D_nE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_E_SI_SDFCHK, nCN_nD_E_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SI_SDFCHK, nCN_nD_nE_SI, 1'b1);
    tsmc_xbuf (CN_D_E_nSI_SDFCHK, CN_D_E_nSI, 1'b1);
    tsmc_xbuf (CN_D_nE_nSI_SDFCHK, CN_D_nE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nE_nSI_SDFCHK, CN_nD_nE_nSI, 1'b1);
    tsmc_xbuf (CN_D_E_SE_SDFCHK, CN_D_E_SE, 1'b1);
    tsmc_xbuf (CN_D_nE_SE_SDFCHK, CN_D_nE_SE, 1'b1);
    tsmc_xbuf (CN_nD_nE_SE_SDFCHK, CN_nD_nE_SE, 1'b1);
    tsmc_xbuf (CN_nD_E_SE_SDFCHK, CN_nD_E_SE, 1'b1);
    tsmc_xbuf (nCN_D_E_SE_SDFCHK, nCN_D_E_SE, 1'b1);
    tsmc_xbuf (nCN_D_nE_SE_SDFCHK, nCN_D_nE_SE, 1'b1);
    tsmc_xbuf (nCN_nD_E_SE_SDFCHK, nCN_nD_E_SE, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SE_SDFCHK, nCN_nD_nE_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    not (nE, E);
    and (CN_D_E_SE_SI, CN, D, E, SE, SI);
    and (CN_D_E_nSE_SI, CN, D, E, nSE, SI);
    and (CN_D_E_nSE_nSI, CN, D, E, nSE, nSI);
    and (CN_nD_E_SE_SI, CN, nD, E, SE, SI);
    and (nCN_D_E_SE_SI, nCN, D, E, SE, SI);
    and (nCN_D_nE_SE_SI, nCN, D, nE, SE, SI);
    and (nCN_nD_E_SE_SI, nCN, nD, E, SE, SI);
    and (nCN_nD_nE_SE_SI, nCN, nD, nE, SE, SI);
    and (CN_D_nE_SE_SI, CN, D, nE, SE, SI);
    and (CN_nD_nE_SE_SI, CN, nD, nE, SE, SI);
    and (CN_D_E_SE_nSI, CN, D, E, SE, nSI);
    and (CN_nD_E_SE_nSI, CN, nD, E, SE, nSI);
    and (CN_nD_E_nSE_SI, CN, nD, E, nSE, SI);
    and (CN_nD_E_nSE_nSI, CN, nD, E, nSE, nSI);
    and (nCN_D_E_SE_nSI, nCN, D, E, SE, nSI);
    and (nCN_D_E_nSE_SI, nCN, D, E, nSE, SI);
    and (nCN_D_E_nSE_nSI, nCN, D, E, nSE, nSI);
    and (nCN_D_nE_SE_nSI, nCN, D, nE, SE, nSI);
    and (nCN_D_nE_nSE_SI, nCN, D, nE, nSE, SI);
    and (nCN_D_nE_nSE_nSI, nCN, D, nE, nSE, nSI);
    and (nCN_nD_E_SE_nSI, nCN, nD, E, SE, nSI);
    and (nCN_nD_E_nSE_SI, nCN, nD, E, nSE, SI);
    and (nCN_nD_E_nSE_nSI, nCN, nD, E, nSE, nSI);
    and (nCN_nD_nE_SE_nSI, nCN, nD, nE, SE, nSI);
    and (nCN_nD_nE_nSE_SI, nCN, nD, nE, nSE, SI);
    and (nCN_nD_nE_nSE_nSI, nCN, nD, nE, nSE, nSI);
    and (CN_D_nE_SE_nSI, CN, D, nE, SE, nSI);
    and (CN_nD_nE_SE_nSI, CN, nD, nE, SE, nSI);
    and (D_E_nSE_SI, D, E, nSE, SI);
    and (D_E_nSE_nSI, D, E, nSE, nSI);
    and (D_nE_nSE_SI, D, nE, nSE, SI);
    and (D_nE_nSE_nSI, D, nE, nSE, nSI);
    and (nD_nE_nSE_SI, nD, nE, nSE, SI);
    and (nD_nE_nSE_nSI, nD, nE, nSE, nSI);
    and (CN_E_nSE_SI, CN, E, nSE, SI);
    and (CN_E_nSE_nSI, CN, E, nSE, nSI);
    and (CN_D_nSE_SI, CN, D, nSE, SI);
    and (CN_D_nSE_nSI, CN, D, nSE, nSI);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);
    and (CN_D_nE_SI, CN, D, nE, SI);
    and (CN_nD_nE_SI, CN, nD, nE, SI);
    and (CN_nD_E_SI, CN, nD, E, SI);
    and (nCN_D_E_SI, nCN, D, E, SI);
    and (nCN_D_nE_SI, nCN, D, nE, SI);
    and (nCN_nD_E_SI, nCN, nD, E, SI);
    and (nCN_nD_nE_SI, nCN, nD, nE, SI);
    and (CN_D_E_nSI, CN, D, E, nSI);
    and (CN_D_nE_nSI, CN, D, nE, nSI);
    and (CN_nD_nE_nSI, CN, nD, nE, nSI);
    and (CN_D_E_SE, CN, D, E, SE);
    and (CN_D_nE_SE, CN, D, nE, SE);
    and (CN_nD_nE_SE, CN, nD, nE, SE);
    and (CN_nD_E_SE, CN, nD, E, SE);
    and (nCN_D_E_SE, nCN, D, E, SE);
    and (nCN_D_nE_SE, nCN, D, nE, SE);
    and (nCN_nD_E_SE, nCN, nD, E, SE);
    and (nCN_nD_nE_SE, nCN, nD, nE, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    and  (D_check, E_d, CN_d, SE_int_not);
    and  (E_check, CN_d, SE_int_not);
    buf  (SI_check, SE_d);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    and  (D_check, E, CN, SE_int_not);
    and  (E_check, CN, SE_int_not);
    buf  (SI_check, SE);
  `endif
  buf  (CN_check, SE_int_not);
  or   (CP_check, D_check, E_check, CN_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && E && D) || (!(SE) && CN && !(E) && Q_buf)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && CN && E && D) || (!(SE) && CN && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_E_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_E_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_E_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_E_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_E_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFKCND1 (SI, D, E, SE, CP, CN, Q, QN);
    input SI, D, SE, CP, CN, E;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d, E_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        and (D2, CN_d, D1);
        tsmc_mux (D3, D2, SI_d, SE_d);
        tsmc_dff (Q_buf, D3, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        and (D2, CN, D1);
        tsmc_mux (D3, D2, SI, SE);
        tsmc_dff (Q_buf, D3, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_E_SE_SI_SDFCHK, CN_D_E_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_E_nSE_SI_SDFCHK, CN_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (CN_D_E_nSE_nSI_SDFCHK, CN_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_E_SE_SI_SDFCHK, CN_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nCN_D_E_SE_SI_SDFCHK, nCN_D_E_SE_SI, 1'b1);
    tsmc_xbuf (nCN_D_nE_SE_SI_SDFCHK, nCN_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_E_SE_SI_SDFCHK, nCN_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SE_SI_SDFCHK, nCN_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_nE_SE_SI_SDFCHK, CN_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nE_SE_SI_SDFCHK, CN_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_E_SE_nSI_SDFCHK, CN_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_E_SE_nSI_SDFCHK, CN_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_E_nSE_SI_SDFCHK, CN_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_E_nSE_nSI_SDFCHK, CN_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_E_SE_nSI_SDFCHK, nCN_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_E_nSE_SI_SDFCHK, nCN_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_D_E_nSE_nSI_SDFCHK, nCN_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_nE_SE_nSI_SDFCHK, nCN_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_nE_nSE_SI_SDFCHK, nCN_D_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_D_nE_nSE_nSI_SDFCHK, nCN_D_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_E_SE_nSI_SDFCHK, nCN_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_E_nSE_SI_SDFCHK, nCN_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_E_nSE_nSI_SDFCHK, nCN_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SE_nSI_SDFCHK, nCN_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_nSE_SI_SDFCHK, nCN_nD_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_nSE_nSI_SDFCHK, nCN_nD_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_D_nE_SE_nSI_SDFCHK, CN_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nE_SE_nSI_SDFCHK, CN_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (D_E_nSE_SI_SDFCHK, D_E_nSE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_nSI_SDFCHK, D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nE_nSE_SI_SDFCHK, D_nE_nSE_SI, 1'b1);
    tsmc_xbuf (D_nE_nSE_nSI_SDFCHK, D_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_nSE_SI_SDFCHK, nD_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nE_nSE_nSI_SDFCHK, nD_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_E_nSE_SI_SDFCHK, CN_E_nSE_SI, 1'b1);
    tsmc_xbuf (CN_E_nSE_nSI_SDFCHK, CN_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SDFCHK, CN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SDFCHK, CN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_D_nE_SI_SDFCHK, CN_D_nE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nE_SI_SDFCHK, CN_nD_nE_SI, 1'b1);
    tsmc_xbuf (CN_nD_E_SI_SDFCHK, CN_nD_E_SI, 1'b1);
    tsmc_xbuf (nCN_D_E_SI_SDFCHK, nCN_D_E_SI, 1'b1);
    tsmc_xbuf (nCN_D_nE_SI_SDFCHK, nCN_D_nE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_E_SI_SDFCHK, nCN_nD_E_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SI_SDFCHK, nCN_nD_nE_SI, 1'b1);
    tsmc_xbuf (CN_D_E_nSI_SDFCHK, CN_D_E_nSI, 1'b1);
    tsmc_xbuf (CN_D_nE_nSI_SDFCHK, CN_D_nE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nE_nSI_SDFCHK, CN_nD_nE_nSI, 1'b1);
    tsmc_xbuf (CN_D_E_SE_SDFCHK, CN_D_E_SE, 1'b1);
    tsmc_xbuf (CN_nD_E_SE_SDFCHK, CN_nD_E_SE, 1'b1);
    tsmc_xbuf (nCN_D_E_SE_SDFCHK, nCN_D_E_SE, 1'b1);
    tsmc_xbuf (nCN_D_nE_SE_SDFCHK, nCN_D_nE_SE, 1'b1);
    tsmc_xbuf (nCN_nD_E_SE_SDFCHK, nCN_nD_E_SE, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SE_SDFCHK, nCN_nD_nE_SE, 1'b1);
    tsmc_xbuf (CN_D_nE_SE_SDFCHK, CN_D_nE_SE, 1'b1);
    tsmc_xbuf (CN_nD_nE_SE_SDFCHK, CN_nD_nE_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    not (nE, E);
    and (CN_D_E_SE_SI, CN, D, E, SE, SI);
    and (CN_D_E_nSE_SI, CN, D, E, nSE, SI);
    and (CN_D_E_nSE_nSI, CN, D, E, nSE, nSI);
    and (CN_nD_E_SE_SI, CN, nD, E, SE, SI);
    and (nCN_D_E_SE_SI, nCN, D, E, SE, SI);
    and (nCN_D_nE_SE_SI, nCN, D, nE, SE, SI);
    and (nCN_nD_E_SE_SI, nCN, nD, E, SE, SI);
    and (nCN_nD_nE_SE_SI, nCN, nD, nE, SE, SI);
    and (CN_D_nE_SE_SI, CN, D, nE, SE, SI);
    and (CN_nD_nE_SE_SI, CN, nD, nE, SE, SI);
    and (CN_D_E_SE_nSI, CN, D, E, SE, nSI);
    and (CN_nD_E_SE_nSI, CN, nD, E, SE, nSI);
    and (CN_nD_E_nSE_SI, CN, nD, E, nSE, SI);
    and (CN_nD_E_nSE_nSI, CN, nD, E, nSE, nSI);
    and (nCN_D_E_SE_nSI, nCN, D, E, SE, nSI);
    and (nCN_D_E_nSE_SI, nCN, D, E, nSE, SI);
    and (nCN_D_E_nSE_nSI, nCN, D, E, nSE, nSI);
    and (nCN_D_nE_SE_nSI, nCN, D, nE, SE, nSI);
    and (nCN_D_nE_nSE_SI, nCN, D, nE, nSE, SI);
    and (nCN_D_nE_nSE_nSI, nCN, D, nE, nSE, nSI);
    and (nCN_nD_E_SE_nSI, nCN, nD, E, SE, nSI);
    and (nCN_nD_E_nSE_SI, nCN, nD, E, nSE, SI);
    and (nCN_nD_E_nSE_nSI, nCN, nD, E, nSE, nSI);
    and (nCN_nD_nE_SE_nSI, nCN, nD, nE, SE, nSI);
    and (nCN_nD_nE_nSE_SI, nCN, nD, nE, nSE, SI);
    and (nCN_nD_nE_nSE_nSI, nCN, nD, nE, nSE, nSI);
    and (CN_D_nE_SE_nSI, CN, D, nE, SE, nSI);
    and (CN_nD_nE_SE_nSI, CN, nD, nE, SE, nSI);
    and (D_E_nSE_SI, D, E, nSE, SI);
    and (D_E_nSE_nSI, D, E, nSE, nSI);
    and (D_nE_nSE_SI, D, nE, nSE, SI);
    and (D_nE_nSE_nSI, D, nE, nSE, nSI);
    and (nD_nE_nSE_SI, nD, nE, nSE, SI);
    and (nD_nE_nSE_nSI, nD, nE, nSE, nSI);
    and (CN_E_nSE_SI, CN, E, nSE, SI);
    and (CN_E_nSE_nSI, CN, E, nSE, nSI);
    and (CN_D_nSE_SI, CN, D, nSE, SI);
    and (CN_D_nSE_nSI, CN, D, nSE, nSI);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);
    and (CN_D_nE_SI, CN, D, nE, SI);
    and (CN_nD_nE_SI, CN, nD, nE, SI);
    and (CN_nD_E_SI, CN, nD, E, SI);
    and (nCN_D_E_SI, nCN, D, E, SI);
    and (nCN_D_nE_SI, nCN, D, nE, SI);
    and (nCN_nD_E_SI, nCN, nD, E, SI);
    and (nCN_nD_nE_SI, nCN, nD, nE, SI);
    and (CN_D_E_nSI, CN, D, E, nSI);
    and (CN_D_nE_nSI, CN, D, nE, nSI);
    and (CN_nD_nE_nSI, CN, nD, nE, nSI);
    and (CN_D_E_SE, CN, D, E, SE);
    and (CN_nD_E_SE, CN, nD, E, SE);
    and (nCN_D_E_SE, nCN, D, E, SE);
    and (nCN_D_nE_SE, nCN, D, nE, SE);
    and (nCN_nD_E_SE, nCN, nD, E, SE);
    and (nCN_nD_nE_SE, nCN, nD, nE, SE);
    and (CN_D_nE_SE, CN, D, nE, SE);
    and (CN_nD_nE_SE, CN, nD, nE, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    and  (D_check, E_d, CN_d, SE_int_not);
    and  (E_check, CN_d, SE_int_not);
    buf  (SI_check, SE_d);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    and  (D_check, E, CN, SE_int_not);
    and  (E_check, CN, SE_int_not);
    buf  (SI_check, SE);
  `endif
  buf  (CN_check, SE_int_not);
  or   (CP_check, D_check, E_check, CN_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && E && D) || (!(SE) && CN && !(E) && Q_buf)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && CN && E && D) || (!(SE) && CN && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_E_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_E_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_E_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_E_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_E_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFKCND2 (SI, D, E, SE, CP, CN, Q, QN);
    input SI, D, SE, CP, CN, E;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d, E_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        and (D2, CN_d, D1);
        tsmc_mux (D3, D2, SI_d, SE_d);
        tsmc_dff (Q_buf, D3, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        and (D2, CN, D1);
        tsmc_mux (D3, D2, SI, SE);
        tsmc_dff (Q_buf, D3, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_E_SE_SI_SDFCHK, CN_D_E_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_E_nSE_SI_SDFCHK, CN_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (CN_D_E_nSE_nSI_SDFCHK, CN_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_E_SE_SI_SDFCHK, CN_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nCN_D_E_SE_SI_SDFCHK, nCN_D_E_SE_SI, 1'b1);
    tsmc_xbuf (nCN_D_nE_SE_SI_SDFCHK, nCN_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_E_SE_SI_SDFCHK, nCN_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SE_SI_SDFCHK, nCN_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_nE_SE_SI_SDFCHK, CN_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nE_SE_SI_SDFCHK, CN_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_E_SE_nSI_SDFCHK, CN_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_E_SE_nSI_SDFCHK, CN_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_E_nSE_SI_SDFCHK, CN_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_E_nSE_nSI_SDFCHK, CN_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_E_SE_nSI_SDFCHK, nCN_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_E_nSE_SI_SDFCHK, nCN_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_D_E_nSE_nSI_SDFCHK, nCN_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_nE_SE_nSI_SDFCHK, nCN_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_nE_nSE_SI_SDFCHK, nCN_D_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_D_nE_nSE_nSI_SDFCHK, nCN_D_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_E_SE_nSI_SDFCHK, nCN_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_E_nSE_SI_SDFCHK, nCN_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_E_nSE_nSI_SDFCHK, nCN_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SE_nSI_SDFCHK, nCN_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_nSE_SI_SDFCHK, nCN_nD_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_nSE_nSI_SDFCHK, nCN_nD_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_D_nE_SE_nSI_SDFCHK, CN_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nE_SE_nSI_SDFCHK, CN_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (D_E_nSE_SI_SDFCHK, D_E_nSE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_nSI_SDFCHK, D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nE_nSE_SI_SDFCHK, D_nE_nSE_SI, 1'b1);
    tsmc_xbuf (D_nE_nSE_nSI_SDFCHK, D_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_nSE_SI_SDFCHK, nD_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nE_nSE_nSI_SDFCHK, nD_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_E_nSE_SI_SDFCHK, CN_E_nSE_SI, 1'b1);
    tsmc_xbuf (CN_E_nSE_nSI_SDFCHK, CN_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SDFCHK, CN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SDFCHK, CN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_D_nE_SI_SDFCHK, CN_D_nE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nE_SI_SDFCHK, CN_nD_nE_SI, 1'b1);
    tsmc_xbuf (CN_nD_E_SI_SDFCHK, CN_nD_E_SI, 1'b1);
    tsmc_xbuf (nCN_D_E_SI_SDFCHK, nCN_D_E_SI, 1'b1);
    tsmc_xbuf (nCN_D_nE_SI_SDFCHK, nCN_D_nE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_E_SI_SDFCHK, nCN_nD_E_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SI_SDFCHK, nCN_nD_nE_SI, 1'b1);
    tsmc_xbuf (CN_D_E_nSI_SDFCHK, CN_D_E_nSI, 1'b1);
    tsmc_xbuf (CN_D_nE_nSI_SDFCHK, CN_D_nE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nE_nSI_SDFCHK, CN_nD_nE_nSI, 1'b1);
    tsmc_xbuf (CN_D_E_SE_SDFCHK, CN_D_E_SE, 1'b1);
    tsmc_xbuf (CN_nD_E_SE_SDFCHK, CN_nD_E_SE, 1'b1);
    tsmc_xbuf (nCN_D_E_SE_SDFCHK, nCN_D_E_SE, 1'b1);
    tsmc_xbuf (nCN_D_nE_SE_SDFCHK, nCN_D_nE_SE, 1'b1);
    tsmc_xbuf (nCN_nD_E_SE_SDFCHK, nCN_nD_E_SE, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SE_SDFCHK, nCN_nD_nE_SE, 1'b1);
    tsmc_xbuf (CN_D_nE_SE_SDFCHK, CN_D_nE_SE, 1'b1);
    tsmc_xbuf (CN_nD_nE_SE_SDFCHK, CN_nD_nE_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    not (nE, E);
    and (CN_D_E_SE_SI, CN, D, E, SE, SI);
    and (CN_D_E_nSE_SI, CN, D, E, nSE, SI);
    and (CN_D_E_nSE_nSI, CN, D, E, nSE, nSI);
    and (CN_nD_E_SE_SI, CN, nD, E, SE, SI);
    and (nCN_D_E_SE_SI, nCN, D, E, SE, SI);
    and (nCN_D_nE_SE_SI, nCN, D, nE, SE, SI);
    and (nCN_nD_E_SE_SI, nCN, nD, E, SE, SI);
    and (nCN_nD_nE_SE_SI, nCN, nD, nE, SE, SI);
    and (CN_D_nE_SE_SI, CN, D, nE, SE, SI);
    and (CN_nD_nE_SE_SI, CN, nD, nE, SE, SI);
    and (CN_D_E_SE_nSI, CN, D, E, SE, nSI);
    and (CN_nD_E_SE_nSI, CN, nD, E, SE, nSI);
    and (CN_nD_E_nSE_SI, CN, nD, E, nSE, SI);
    and (CN_nD_E_nSE_nSI, CN, nD, E, nSE, nSI);
    and (nCN_D_E_SE_nSI, nCN, D, E, SE, nSI);
    and (nCN_D_E_nSE_SI, nCN, D, E, nSE, SI);
    and (nCN_D_E_nSE_nSI, nCN, D, E, nSE, nSI);
    and (nCN_D_nE_SE_nSI, nCN, D, nE, SE, nSI);
    and (nCN_D_nE_nSE_SI, nCN, D, nE, nSE, SI);
    and (nCN_D_nE_nSE_nSI, nCN, D, nE, nSE, nSI);
    and (nCN_nD_E_SE_nSI, nCN, nD, E, SE, nSI);
    and (nCN_nD_E_nSE_SI, nCN, nD, E, nSE, SI);
    and (nCN_nD_E_nSE_nSI, nCN, nD, E, nSE, nSI);
    and (nCN_nD_nE_SE_nSI, nCN, nD, nE, SE, nSI);
    and (nCN_nD_nE_nSE_SI, nCN, nD, nE, nSE, SI);
    and (nCN_nD_nE_nSE_nSI, nCN, nD, nE, nSE, nSI);
    and (CN_D_nE_SE_nSI, CN, D, nE, SE, nSI);
    and (CN_nD_nE_SE_nSI, CN, nD, nE, SE, nSI);
    and (D_E_nSE_SI, D, E, nSE, SI);
    and (D_E_nSE_nSI, D, E, nSE, nSI);
    and (D_nE_nSE_SI, D, nE, nSE, SI);
    and (D_nE_nSE_nSI, D, nE, nSE, nSI);
    and (nD_nE_nSE_SI, nD, nE, nSE, SI);
    and (nD_nE_nSE_nSI, nD, nE, nSE, nSI);
    and (CN_E_nSE_SI, CN, E, nSE, SI);
    and (CN_E_nSE_nSI, CN, E, nSE, nSI);
    and (CN_D_nSE_SI, CN, D, nSE, SI);
    and (CN_D_nSE_nSI, CN, D, nSE, nSI);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);
    and (CN_D_nE_SI, CN, D, nE, SI);
    and (CN_nD_nE_SI, CN, nD, nE, SI);
    and (CN_nD_E_SI, CN, nD, E, SI);
    and (nCN_D_E_SI, nCN, D, E, SI);
    and (nCN_D_nE_SI, nCN, D, nE, SI);
    and (nCN_nD_E_SI, nCN, nD, E, SI);
    and (nCN_nD_nE_SI, nCN, nD, nE, SI);
    and (CN_D_E_nSI, CN, D, E, nSI);
    and (CN_D_nE_nSI, CN, D, nE, nSI);
    and (CN_nD_nE_nSI, CN, nD, nE, nSI);
    and (CN_D_E_SE, CN, D, E, SE);
    and (CN_nD_E_SE, CN, nD, E, SE);
    and (nCN_D_E_SE, nCN, D, E, SE);
    and (nCN_D_nE_SE, nCN, D, nE, SE);
    and (nCN_nD_E_SE, nCN, nD, E, SE);
    and (nCN_nD_nE_SE, nCN, nD, nE, SE);
    and (CN_D_nE_SE, CN, D, nE, SE);
    and (CN_nD_nE_SE, CN, nD, nE, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    and  (D_check, E_d, CN_d, SE_int_not);
    and  (E_check, CN_d, SE_int_not);
    buf  (SI_check, SE_d);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    and  (D_check, E, CN, SE_int_not);
    and  (E_check, CN, SE_int_not);
    buf  (SI_check, SE);
  `endif
  buf  (CN_check, SE_int_not);
  or   (CP_check, D_check, E_check, CN_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && E && D) || (!(SE) && CN && !(E) && Q_buf)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && CN && E && D) || (!(SE) && CN && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_E_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_E_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_E_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_E_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_E_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFKCND4 (SI, D, E, SE, CP, CN, Q, QN);
    input SI, D, SE, CP, CN, E;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d, E_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        and (D2, CN_d, D1);
        tsmc_mux (D3, D2, SI_d, SE_d);
        tsmc_dff (Q_buf, D3, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        and (D2, CN, D1);
        tsmc_mux (D3, D2, SI, SE);
        tsmc_dff (Q_buf, D3, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_E_SE_SI_SDFCHK, CN_D_E_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_E_nSE_SI_SDFCHK, CN_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (CN_D_E_nSE_nSI_SDFCHK, CN_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_E_SE_SI_SDFCHK, CN_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nCN_D_E_SE_SI_SDFCHK, nCN_D_E_SE_SI, 1'b1);
    tsmc_xbuf (nCN_D_nE_SE_SI_SDFCHK, nCN_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_E_SE_SI_SDFCHK, nCN_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SE_SI_SDFCHK, nCN_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_nE_SE_SI_SDFCHK, CN_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nE_SE_SI_SDFCHK, CN_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_E_SE_nSI_SDFCHK, CN_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_E_SE_nSI_SDFCHK, CN_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_E_nSE_SI_SDFCHK, CN_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_E_nSE_nSI_SDFCHK, CN_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_E_SE_nSI_SDFCHK, nCN_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_E_nSE_SI_SDFCHK, nCN_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_D_E_nSE_nSI_SDFCHK, nCN_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_nE_SE_nSI_SDFCHK, nCN_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_nE_nSE_SI_SDFCHK, nCN_D_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_D_nE_nSE_nSI_SDFCHK, nCN_D_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_E_SE_nSI_SDFCHK, nCN_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_E_nSE_SI_SDFCHK, nCN_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_E_nSE_nSI_SDFCHK, nCN_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SE_nSI_SDFCHK, nCN_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_nSE_SI_SDFCHK, nCN_nD_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_nSE_nSI_SDFCHK, nCN_nD_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_D_nE_SE_nSI_SDFCHK, CN_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nE_SE_nSI_SDFCHK, CN_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (D_E_nSE_SI_SDFCHK, D_E_nSE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_nSI_SDFCHK, D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nE_nSE_SI_SDFCHK, D_nE_nSE_SI, 1'b1);
    tsmc_xbuf (D_nE_nSE_nSI_SDFCHK, D_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_nSE_SI_SDFCHK, nD_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nE_nSE_nSI_SDFCHK, nD_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_E_nSE_SI_SDFCHK, CN_E_nSE_SI, 1'b1);
    tsmc_xbuf (CN_E_nSE_nSI_SDFCHK, CN_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SDFCHK, CN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SDFCHK, CN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_D_nE_SI_SDFCHK, CN_D_nE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nE_SI_SDFCHK, CN_nD_nE_SI, 1'b1);
    tsmc_xbuf (CN_nD_E_SI_SDFCHK, CN_nD_E_SI, 1'b1);
    tsmc_xbuf (nCN_D_E_SI_SDFCHK, nCN_D_E_SI, 1'b1);
    tsmc_xbuf (nCN_D_nE_SI_SDFCHK, nCN_D_nE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_E_SI_SDFCHK, nCN_nD_E_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SI_SDFCHK, nCN_nD_nE_SI, 1'b1);
    tsmc_xbuf (CN_D_E_nSI_SDFCHK, CN_D_E_nSI, 1'b1);
    tsmc_xbuf (CN_D_nE_nSI_SDFCHK, CN_D_nE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nE_nSI_SDFCHK, CN_nD_nE_nSI, 1'b1);
    tsmc_xbuf (CN_D_E_SE_SDFCHK, CN_D_E_SE, 1'b1);
    tsmc_xbuf (CN_nD_E_SE_SDFCHK, CN_nD_E_SE, 1'b1);
    tsmc_xbuf (nCN_D_E_SE_SDFCHK, nCN_D_E_SE, 1'b1);
    tsmc_xbuf (nCN_D_nE_SE_SDFCHK, nCN_D_nE_SE, 1'b1);
    tsmc_xbuf (nCN_nD_E_SE_SDFCHK, nCN_nD_E_SE, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SE_SDFCHK, nCN_nD_nE_SE, 1'b1);
    tsmc_xbuf (CN_D_nE_SE_SDFCHK, CN_D_nE_SE, 1'b1);
    tsmc_xbuf (CN_nD_nE_SE_SDFCHK, CN_nD_nE_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    not (nE, E);
    and (CN_D_E_SE_SI, CN, D, E, SE, SI);
    and (CN_D_E_nSE_SI, CN, D, E, nSE, SI);
    and (CN_D_E_nSE_nSI, CN, D, E, nSE, nSI);
    and (CN_nD_E_SE_SI, CN, nD, E, SE, SI);
    and (nCN_D_E_SE_SI, nCN, D, E, SE, SI);
    and (nCN_D_nE_SE_SI, nCN, D, nE, SE, SI);
    and (nCN_nD_E_SE_SI, nCN, nD, E, SE, SI);
    and (nCN_nD_nE_SE_SI, nCN, nD, nE, SE, SI);
    and (CN_D_nE_SE_SI, CN, D, nE, SE, SI);
    and (CN_nD_nE_SE_SI, CN, nD, nE, SE, SI);
    and (CN_D_E_SE_nSI, CN, D, E, SE, nSI);
    and (CN_nD_E_SE_nSI, CN, nD, E, SE, nSI);
    and (CN_nD_E_nSE_SI, CN, nD, E, nSE, SI);
    and (CN_nD_E_nSE_nSI, CN, nD, E, nSE, nSI);
    and (nCN_D_E_SE_nSI, nCN, D, E, SE, nSI);
    and (nCN_D_E_nSE_SI, nCN, D, E, nSE, SI);
    and (nCN_D_E_nSE_nSI, nCN, D, E, nSE, nSI);
    and (nCN_D_nE_SE_nSI, nCN, D, nE, SE, nSI);
    and (nCN_D_nE_nSE_SI, nCN, D, nE, nSE, SI);
    and (nCN_D_nE_nSE_nSI, nCN, D, nE, nSE, nSI);
    and (nCN_nD_E_SE_nSI, nCN, nD, E, SE, nSI);
    and (nCN_nD_E_nSE_SI, nCN, nD, E, nSE, SI);
    and (nCN_nD_E_nSE_nSI, nCN, nD, E, nSE, nSI);
    and (nCN_nD_nE_SE_nSI, nCN, nD, nE, SE, nSI);
    and (nCN_nD_nE_nSE_SI, nCN, nD, nE, nSE, SI);
    and (nCN_nD_nE_nSE_nSI, nCN, nD, nE, nSE, nSI);
    and (CN_D_nE_SE_nSI, CN, D, nE, SE, nSI);
    and (CN_nD_nE_SE_nSI, CN, nD, nE, SE, nSI);
    and (D_E_nSE_SI, D, E, nSE, SI);
    and (D_E_nSE_nSI, D, E, nSE, nSI);
    and (D_nE_nSE_SI, D, nE, nSE, SI);
    and (D_nE_nSE_nSI, D, nE, nSE, nSI);
    and (nD_nE_nSE_SI, nD, nE, nSE, SI);
    and (nD_nE_nSE_nSI, nD, nE, nSE, nSI);
    and (CN_E_nSE_SI, CN, E, nSE, SI);
    and (CN_E_nSE_nSI, CN, E, nSE, nSI);
    and (CN_D_nSE_SI, CN, D, nSE, SI);
    and (CN_D_nSE_nSI, CN, D, nSE, nSI);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);
    and (CN_D_nE_SI, CN, D, nE, SI);
    and (CN_nD_nE_SI, CN, nD, nE, SI);
    and (CN_nD_E_SI, CN, nD, E, SI);
    and (nCN_D_E_SI, nCN, D, E, SI);
    and (nCN_D_nE_SI, nCN, D, nE, SI);
    and (nCN_nD_E_SI, nCN, nD, E, SI);
    and (nCN_nD_nE_SI, nCN, nD, nE, SI);
    and (CN_D_E_nSI, CN, D, E, nSI);
    and (CN_D_nE_nSI, CN, D, nE, nSI);
    and (CN_nD_nE_nSI, CN, nD, nE, nSI);
    and (CN_D_E_SE, CN, D, E, SE);
    and (CN_nD_E_SE, CN, nD, E, SE);
    and (nCN_D_E_SE, nCN, D, E, SE);
    and (nCN_D_nE_SE, nCN, D, nE, SE);
    and (nCN_nD_E_SE, nCN, nD, E, SE);
    and (nCN_nD_nE_SE, nCN, nD, nE, SE);
    and (CN_D_nE_SE, CN, D, nE, SE);
    and (CN_nD_nE_SE, CN, nD, nE, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    and  (D_check, E_d, CN_d, SE_int_not);
    and  (E_check, CN_d, SE_int_not);
    buf  (SI_check, SE_d);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    and  (D_check, E, CN, SE_int_not);
    and  (E_check, CN, SE_int_not);
    buf  (SI_check, SE);
  `endif
  buf  (CN_check, SE_int_not);
  or   (CP_check, D_check, E_check, CN_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && E && D) || (!(SE) && CN && !(E) && Q_buf)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && CN && E && D) || (!(SE) && CN && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_E_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_E_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_E_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_E_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_E_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFKCNQD0 (SI, D, E, SE, CP, CN, Q);
    input SI, D, SE, CP, CN, E;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d, E_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        and (D2, CN_d, D1);
        tsmc_mux (D3, D2, SI_d, SE_d);
        tsmc_dff (Q_buf, D3, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        and (D2, CN, D1);
        tsmc_mux (D3, D2, SI, SE);
        tsmc_dff (Q_buf, D3, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_E_SE_SI_SDFCHK, CN_D_E_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_E_nSE_SI_SDFCHK, CN_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (CN_D_E_nSE_nSI_SDFCHK, CN_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_E_SE_SI_SDFCHK, CN_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nCN_D_E_SE_SI_SDFCHK, nCN_D_E_SE_SI, 1'b1);
    tsmc_xbuf (nCN_D_nE_SE_SI_SDFCHK, nCN_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_E_SE_SI_SDFCHK, nCN_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SE_SI_SDFCHK, nCN_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_nE_SE_SI_SDFCHK, CN_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nE_SE_SI_SDFCHK, CN_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_E_SE_nSI_SDFCHK, CN_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_E_SE_nSI_SDFCHK, CN_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_E_nSE_SI_SDFCHK, CN_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_E_nSE_nSI_SDFCHK, CN_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_E_SE_nSI_SDFCHK, nCN_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_E_nSE_SI_SDFCHK, nCN_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_D_E_nSE_nSI_SDFCHK, nCN_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_nE_SE_nSI_SDFCHK, nCN_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_nE_nSE_SI_SDFCHK, nCN_D_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_D_nE_nSE_nSI_SDFCHK, nCN_D_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_E_SE_nSI_SDFCHK, nCN_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_E_nSE_SI_SDFCHK, nCN_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_E_nSE_nSI_SDFCHK, nCN_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SE_nSI_SDFCHK, nCN_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_nSE_SI_SDFCHK, nCN_nD_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_nSE_nSI_SDFCHK, nCN_nD_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_D_nE_SE_nSI_SDFCHK, CN_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nE_SE_nSI_SDFCHK, CN_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (D_E_nSE_SI_SDFCHK, D_E_nSE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_nSI_SDFCHK, D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nE_nSE_SI_SDFCHK, D_nE_nSE_SI, 1'b1);
    tsmc_xbuf (D_nE_nSE_nSI_SDFCHK, D_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_nSE_SI_SDFCHK, nD_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nE_nSE_nSI_SDFCHK, nD_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_E_nSE_SI_SDFCHK, CN_E_nSE_SI, 1'b1);
    tsmc_xbuf (CN_E_nSE_nSI_SDFCHK, CN_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SDFCHK, CN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SDFCHK, CN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_D_nE_SI_SDFCHK, CN_D_nE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nE_SI_SDFCHK, CN_nD_nE_SI, 1'b1);
    tsmc_xbuf (CN_nD_E_SI_SDFCHK, CN_nD_E_SI, 1'b1);
    tsmc_xbuf (nCN_D_E_SI_SDFCHK, nCN_D_E_SI, 1'b1);
    tsmc_xbuf (nCN_D_nE_SI_SDFCHK, nCN_D_nE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_E_SI_SDFCHK, nCN_nD_E_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SI_SDFCHK, nCN_nD_nE_SI, 1'b1);
    tsmc_xbuf (CN_D_E_nSI_SDFCHK, CN_D_E_nSI, 1'b1);
    tsmc_xbuf (CN_D_nE_nSI_SDFCHK, CN_D_nE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nE_nSI_SDFCHK, CN_nD_nE_nSI, 1'b1);
    tsmc_xbuf (CN_D_E_SE_SDFCHK, CN_D_E_SE, 1'b1);
    tsmc_xbuf (CN_D_nE_SE_SDFCHK, CN_D_nE_SE, 1'b1);
    tsmc_xbuf (CN_nD_nE_SE_SDFCHK, CN_nD_nE_SE, 1'b1);
    tsmc_xbuf (CN_nD_E_SE_SDFCHK, CN_nD_E_SE, 1'b1);
    tsmc_xbuf (nCN_D_E_SE_SDFCHK, nCN_D_E_SE, 1'b1);
    tsmc_xbuf (nCN_D_nE_SE_SDFCHK, nCN_D_nE_SE, 1'b1);
    tsmc_xbuf (nCN_nD_E_SE_SDFCHK, nCN_nD_E_SE, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SE_SDFCHK, nCN_nD_nE_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    not (nE, E);
    and (CN_D_E_SE_SI, CN, D, E, SE, SI);
    and (CN_D_E_nSE_SI, CN, D, E, nSE, SI);
    and (CN_D_E_nSE_nSI, CN, D, E, nSE, nSI);
    and (CN_nD_E_SE_SI, CN, nD, E, SE, SI);
    and (nCN_D_E_SE_SI, nCN, D, E, SE, SI);
    and (nCN_D_nE_SE_SI, nCN, D, nE, SE, SI);
    and (nCN_nD_E_SE_SI, nCN, nD, E, SE, SI);
    and (nCN_nD_nE_SE_SI, nCN, nD, nE, SE, SI);
    and (CN_D_nE_SE_SI, CN, D, nE, SE, SI);
    and (CN_nD_nE_SE_SI, CN, nD, nE, SE, SI);
    and (CN_D_E_SE_nSI, CN, D, E, SE, nSI);
    and (CN_nD_E_SE_nSI, CN, nD, E, SE, nSI);
    and (CN_nD_E_nSE_SI, CN, nD, E, nSE, SI);
    and (CN_nD_E_nSE_nSI, CN, nD, E, nSE, nSI);
    and (nCN_D_E_SE_nSI, nCN, D, E, SE, nSI);
    and (nCN_D_E_nSE_SI, nCN, D, E, nSE, SI);
    and (nCN_D_E_nSE_nSI, nCN, D, E, nSE, nSI);
    and (nCN_D_nE_SE_nSI, nCN, D, nE, SE, nSI);
    and (nCN_D_nE_nSE_SI, nCN, D, nE, nSE, SI);
    and (nCN_D_nE_nSE_nSI, nCN, D, nE, nSE, nSI);
    and (nCN_nD_E_SE_nSI, nCN, nD, E, SE, nSI);
    and (nCN_nD_E_nSE_SI, nCN, nD, E, nSE, SI);
    and (nCN_nD_E_nSE_nSI, nCN, nD, E, nSE, nSI);
    and (nCN_nD_nE_SE_nSI, nCN, nD, nE, SE, nSI);
    and (nCN_nD_nE_nSE_SI, nCN, nD, nE, nSE, SI);
    and (nCN_nD_nE_nSE_nSI, nCN, nD, nE, nSE, nSI);
    and (CN_D_nE_SE_nSI, CN, D, nE, SE, nSI);
    and (CN_nD_nE_SE_nSI, CN, nD, nE, SE, nSI);
    and (D_E_nSE_SI, D, E, nSE, SI);
    and (D_E_nSE_nSI, D, E, nSE, nSI);
    and (D_nE_nSE_SI, D, nE, nSE, SI);
    and (D_nE_nSE_nSI, D, nE, nSE, nSI);
    and (nD_nE_nSE_SI, nD, nE, nSE, SI);
    and (nD_nE_nSE_nSI, nD, nE, nSE, nSI);
    and (CN_E_nSE_SI, CN, E, nSE, SI);
    and (CN_E_nSE_nSI, CN, E, nSE, nSI);
    and (CN_D_nSE_SI, CN, D, nSE, SI);
    and (CN_D_nSE_nSI, CN, D, nSE, nSI);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);
    and (CN_D_nE_SI, CN, D, nE, SI);
    and (CN_nD_nE_SI, CN, nD, nE, SI);
    and (CN_nD_E_SI, CN, nD, E, SI);
    and (nCN_D_E_SI, nCN, D, E, SI);
    and (nCN_D_nE_SI, nCN, D, nE, SI);
    and (nCN_nD_E_SI, nCN, nD, E, SI);
    and (nCN_nD_nE_SI, nCN, nD, nE, SI);
    and (CN_D_E_nSI, CN, D, E, nSI);
    and (CN_D_nE_nSI, CN, D, nE, nSI);
    and (CN_nD_nE_nSI, CN, nD, nE, nSI);
    and (CN_D_E_SE, CN, D, E, SE);
    and (CN_D_nE_SE, CN, D, nE, SE);
    and (CN_nD_nE_SE, CN, nD, nE, SE);
    and (CN_nD_E_SE, CN, nD, E, SE);
    and (nCN_D_E_SE, nCN, D, E, SE);
    and (nCN_D_nE_SE, nCN, D, nE, SE);
    and (nCN_nD_E_SE, nCN, nD, E, SE);
    and (nCN_nD_nE_SE, nCN, nD, nE, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    and  (D_check, E_d, CN_d, SE_int_not);
    and  (E_check, CN_d, SE_int_not);
    buf  (SI_check, SE_d);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    and  (D_check, E, CN, SE_int_not);
    and  (E_check, CN, SE_int_not);
    buf  (SI_check, SE);
  `endif
  buf  (CN_check, SE_int_not);
  or   (CP_check, D_check, E_check, CN_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && E && D) || (!(SE) && CN && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_E_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_E_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_E_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_E_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_E_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFKCNQD1 (SI, D, E, SE, CP, CN, Q);
    input SI, D, SE, CP, CN, E;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d, E_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        and (D2, CN_d, D1);
        tsmc_mux (D3, D2, SI_d, SE_d);
        tsmc_dff (Q_buf, D3, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        and (D2, CN, D1);
        tsmc_mux (D3, D2, SI, SE);
        tsmc_dff (Q_buf, D3, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_E_SE_SI_SDFCHK, CN_D_E_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_E_nSE_SI_SDFCHK, CN_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (CN_D_E_nSE_nSI_SDFCHK, CN_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_E_SE_SI_SDFCHK, CN_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nCN_D_E_SE_SI_SDFCHK, nCN_D_E_SE_SI, 1'b1);
    tsmc_xbuf (nCN_D_nE_SE_SI_SDFCHK, nCN_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_E_SE_SI_SDFCHK, nCN_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SE_SI_SDFCHK, nCN_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_nE_SE_SI_SDFCHK, CN_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nE_SE_SI_SDFCHK, CN_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_E_SE_nSI_SDFCHK, CN_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_E_SE_nSI_SDFCHK, CN_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_E_nSE_SI_SDFCHK, CN_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_E_nSE_nSI_SDFCHK, CN_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_E_SE_nSI_SDFCHK, nCN_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_E_nSE_SI_SDFCHK, nCN_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_D_E_nSE_nSI_SDFCHK, nCN_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_nE_SE_nSI_SDFCHK, nCN_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_nE_nSE_SI_SDFCHK, nCN_D_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_D_nE_nSE_nSI_SDFCHK, nCN_D_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_E_SE_nSI_SDFCHK, nCN_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_E_nSE_SI_SDFCHK, nCN_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_E_nSE_nSI_SDFCHK, nCN_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SE_nSI_SDFCHK, nCN_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_nSE_SI_SDFCHK, nCN_nD_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_nSE_nSI_SDFCHK, nCN_nD_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_D_nE_SE_nSI_SDFCHK, CN_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nE_SE_nSI_SDFCHK, CN_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (D_E_nSE_SI_SDFCHK, D_E_nSE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_nSI_SDFCHK, D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nE_nSE_SI_SDFCHK, D_nE_nSE_SI, 1'b1);
    tsmc_xbuf (D_nE_nSE_nSI_SDFCHK, D_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_nSE_SI_SDFCHK, nD_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nE_nSE_nSI_SDFCHK, nD_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_E_nSE_SI_SDFCHK, CN_E_nSE_SI, 1'b1);
    tsmc_xbuf (CN_E_nSE_nSI_SDFCHK, CN_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SDFCHK, CN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SDFCHK, CN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_D_nE_SI_SDFCHK, CN_D_nE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nE_SI_SDFCHK, CN_nD_nE_SI, 1'b1);
    tsmc_xbuf (CN_nD_E_SI_SDFCHK, CN_nD_E_SI, 1'b1);
    tsmc_xbuf (nCN_D_E_SI_SDFCHK, nCN_D_E_SI, 1'b1);
    tsmc_xbuf (nCN_D_nE_SI_SDFCHK, nCN_D_nE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_E_SI_SDFCHK, nCN_nD_E_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SI_SDFCHK, nCN_nD_nE_SI, 1'b1);
    tsmc_xbuf (CN_D_E_nSI_SDFCHK, CN_D_E_nSI, 1'b1);
    tsmc_xbuf (CN_D_nE_nSI_SDFCHK, CN_D_nE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nE_nSI_SDFCHK, CN_nD_nE_nSI, 1'b1);
    tsmc_xbuf (CN_D_E_SE_SDFCHK, CN_D_E_SE, 1'b1);
    tsmc_xbuf (CN_nD_E_SE_SDFCHK, CN_nD_E_SE, 1'b1);
    tsmc_xbuf (nCN_D_E_SE_SDFCHK, nCN_D_E_SE, 1'b1);
    tsmc_xbuf (nCN_D_nE_SE_SDFCHK, nCN_D_nE_SE, 1'b1);
    tsmc_xbuf (nCN_nD_E_SE_SDFCHK, nCN_nD_E_SE, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SE_SDFCHK, nCN_nD_nE_SE, 1'b1);
    tsmc_xbuf (CN_D_nE_SE_SDFCHK, CN_D_nE_SE, 1'b1);
    tsmc_xbuf (CN_nD_nE_SE_SDFCHK, CN_nD_nE_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    not (nE, E);
    and (CN_D_E_SE_SI, CN, D, E, SE, SI);
    and (CN_D_E_nSE_SI, CN, D, E, nSE, SI);
    and (CN_D_E_nSE_nSI, CN, D, E, nSE, nSI);
    and (CN_nD_E_SE_SI, CN, nD, E, SE, SI);
    and (nCN_D_E_SE_SI, nCN, D, E, SE, SI);
    and (nCN_D_nE_SE_SI, nCN, D, nE, SE, SI);
    and (nCN_nD_E_SE_SI, nCN, nD, E, SE, SI);
    and (nCN_nD_nE_SE_SI, nCN, nD, nE, SE, SI);
    and (CN_D_nE_SE_SI, CN, D, nE, SE, SI);
    and (CN_nD_nE_SE_SI, CN, nD, nE, SE, SI);
    and (CN_D_E_SE_nSI, CN, D, E, SE, nSI);
    and (CN_nD_E_SE_nSI, CN, nD, E, SE, nSI);
    and (CN_nD_E_nSE_SI, CN, nD, E, nSE, SI);
    and (CN_nD_E_nSE_nSI, CN, nD, E, nSE, nSI);
    and (nCN_D_E_SE_nSI, nCN, D, E, SE, nSI);
    and (nCN_D_E_nSE_SI, nCN, D, E, nSE, SI);
    and (nCN_D_E_nSE_nSI, nCN, D, E, nSE, nSI);
    and (nCN_D_nE_SE_nSI, nCN, D, nE, SE, nSI);
    and (nCN_D_nE_nSE_SI, nCN, D, nE, nSE, SI);
    and (nCN_D_nE_nSE_nSI, nCN, D, nE, nSE, nSI);
    and (nCN_nD_E_SE_nSI, nCN, nD, E, SE, nSI);
    and (nCN_nD_E_nSE_SI, nCN, nD, E, nSE, SI);
    and (nCN_nD_E_nSE_nSI, nCN, nD, E, nSE, nSI);
    and (nCN_nD_nE_SE_nSI, nCN, nD, nE, SE, nSI);
    and (nCN_nD_nE_nSE_SI, nCN, nD, nE, nSE, SI);
    and (nCN_nD_nE_nSE_nSI, nCN, nD, nE, nSE, nSI);
    and (CN_D_nE_SE_nSI, CN, D, nE, SE, nSI);
    and (CN_nD_nE_SE_nSI, CN, nD, nE, SE, nSI);
    and (D_E_nSE_SI, D, E, nSE, SI);
    and (D_E_nSE_nSI, D, E, nSE, nSI);
    and (D_nE_nSE_SI, D, nE, nSE, SI);
    and (D_nE_nSE_nSI, D, nE, nSE, nSI);
    and (nD_nE_nSE_SI, nD, nE, nSE, SI);
    and (nD_nE_nSE_nSI, nD, nE, nSE, nSI);
    and (CN_E_nSE_SI, CN, E, nSE, SI);
    and (CN_E_nSE_nSI, CN, E, nSE, nSI);
    and (CN_D_nSE_SI, CN, D, nSE, SI);
    and (CN_D_nSE_nSI, CN, D, nSE, nSI);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);
    and (CN_D_nE_SI, CN, D, nE, SI);
    and (CN_nD_nE_SI, CN, nD, nE, SI);
    and (CN_nD_E_SI, CN, nD, E, SI);
    and (nCN_D_E_SI, nCN, D, E, SI);
    and (nCN_D_nE_SI, nCN, D, nE, SI);
    and (nCN_nD_E_SI, nCN, nD, E, SI);
    and (nCN_nD_nE_SI, nCN, nD, nE, SI);
    and (CN_D_E_nSI, CN, D, E, nSI);
    and (CN_D_nE_nSI, CN, D, nE, nSI);
    and (CN_nD_nE_nSI, CN, nD, nE, nSI);
    and (CN_D_E_SE, CN, D, E, SE);
    and (CN_nD_E_SE, CN, nD, E, SE);
    and (nCN_D_E_SE, nCN, D, E, SE);
    and (nCN_D_nE_SE, nCN, D, nE, SE);
    and (nCN_nD_E_SE, nCN, nD, E, SE);
    and (nCN_nD_nE_SE, nCN, nD, nE, SE);
    and (CN_D_nE_SE, CN, D, nE, SE);
    and (CN_nD_nE_SE, CN, nD, nE, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    and  (D_check, E_d, CN_d, SE_int_not);
    and  (E_check, CN_d, SE_int_not);
    buf  (SI_check, SE_d);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    and  (D_check, E, CN, SE_int_not);
    and  (E_check, CN, SE_int_not);
    buf  (SI_check, SE);
  `endif
  buf  (CN_check, SE_int_not);
  or   (CP_check, D_check, E_check, CN_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && E && D) || (!(SE) && CN && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_E_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_E_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_E_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_E_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_E_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFKCNQD2 (SI, D, E, SE, CP, CN, Q);
    input SI, D, SE, CP, CN, E;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d, E_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        and (D2, CN_d, D1);
        tsmc_mux (D3, D2, SI_d, SE_d);
        tsmc_dff (Q_buf, D3, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        and (D2, CN, D1);
        tsmc_mux (D3, D2, SI, SE);
        tsmc_dff (Q_buf, D3, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_E_SE_SI_SDFCHK, CN_D_E_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_E_nSE_SI_SDFCHK, CN_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (CN_D_E_nSE_nSI_SDFCHK, CN_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_E_SE_SI_SDFCHK, CN_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nCN_D_E_SE_SI_SDFCHK, nCN_D_E_SE_SI, 1'b1);
    tsmc_xbuf (nCN_D_nE_SE_SI_SDFCHK, nCN_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_E_SE_SI_SDFCHK, nCN_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SE_SI_SDFCHK, nCN_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_nE_SE_SI_SDFCHK, CN_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nE_SE_SI_SDFCHK, CN_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_E_SE_nSI_SDFCHK, CN_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_E_SE_nSI_SDFCHK, CN_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_E_nSE_SI_SDFCHK, CN_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_E_nSE_nSI_SDFCHK, CN_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_E_SE_nSI_SDFCHK, nCN_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_E_nSE_SI_SDFCHK, nCN_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_D_E_nSE_nSI_SDFCHK, nCN_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_nE_SE_nSI_SDFCHK, nCN_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_nE_nSE_SI_SDFCHK, nCN_D_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_D_nE_nSE_nSI_SDFCHK, nCN_D_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_E_SE_nSI_SDFCHK, nCN_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_E_nSE_SI_SDFCHK, nCN_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_E_nSE_nSI_SDFCHK, nCN_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SE_nSI_SDFCHK, nCN_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_nSE_SI_SDFCHK, nCN_nD_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_nSE_nSI_SDFCHK, nCN_nD_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_D_nE_SE_nSI_SDFCHK, CN_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nE_SE_nSI_SDFCHK, CN_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (D_E_nSE_SI_SDFCHK, D_E_nSE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_nSI_SDFCHK, D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nE_nSE_SI_SDFCHK, D_nE_nSE_SI, 1'b1);
    tsmc_xbuf (D_nE_nSE_nSI_SDFCHK, D_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_nSE_SI_SDFCHK, nD_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nE_nSE_nSI_SDFCHK, nD_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_E_nSE_SI_SDFCHK, CN_E_nSE_SI, 1'b1);
    tsmc_xbuf (CN_E_nSE_nSI_SDFCHK, CN_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SDFCHK, CN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SDFCHK, CN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_D_nE_SI_SDFCHK, CN_D_nE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nE_SI_SDFCHK, CN_nD_nE_SI, 1'b1);
    tsmc_xbuf (CN_nD_E_SI_SDFCHK, CN_nD_E_SI, 1'b1);
    tsmc_xbuf (nCN_D_E_SI_SDFCHK, nCN_D_E_SI, 1'b1);
    tsmc_xbuf (nCN_D_nE_SI_SDFCHK, nCN_D_nE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_E_SI_SDFCHK, nCN_nD_E_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SI_SDFCHK, nCN_nD_nE_SI, 1'b1);
    tsmc_xbuf (CN_D_E_nSI_SDFCHK, CN_D_E_nSI, 1'b1);
    tsmc_xbuf (CN_D_nE_nSI_SDFCHK, CN_D_nE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nE_nSI_SDFCHK, CN_nD_nE_nSI, 1'b1);
    tsmc_xbuf (CN_D_E_SE_SDFCHK, CN_D_E_SE, 1'b1);
    tsmc_xbuf (CN_nD_E_SE_SDFCHK, CN_nD_E_SE, 1'b1);
    tsmc_xbuf (nCN_D_E_SE_SDFCHK, nCN_D_E_SE, 1'b1);
    tsmc_xbuf (nCN_D_nE_SE_SDFCHK, nCN_D_nE_SE, 1'b1);
    tsmc_xbuf (nCN_nD_E_SE_SDFCHK, nCN_nD_E_SE, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SE_SDFCHK, nCN_nD_nE_SE, 1'b1);
    tsmc_xbuf (CN_D_nE_SE_SDFCHK, CN_D_nE_SE, 1'b1);
    tsmc_xbuf (CN_nD_nE_SE_SDFCHK, CN_nD_nE_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    not (nE, E);
    and (CN_D_E_SE_SI, CN, D, E, SE, SI);
    and (CN_D_E_nSE_SI, CN, D, E, nSE, SI);
    and (CN_D_E_nSE_nSI, CN, D, E, nSE, nSI);
    and (CN_nD_E_SE_SI, CN, nD, E, SE, SI);
    and (nCN_D_E_SE_SI, nCN, D, E, SE, SI);
    and (nCN_D_nE_SE_SI, nCN, D, nE, SE, SI);
    and (nCN_nD_E_SE_SI, nCN, nD, E, SE, SI);
    and (nCN_nD_nE_SE_SI, nCN, nD, nE, SE, SI);
    and (CN_D_nE_SE_SI, CN, D, nE, SE, SI);
    and (CN_nD_nE_SE_SI, CN, nD, nE, SE, SI);
    and (CN_D_E_SE_nSI, CN, D, E, SE, nSI);
    and (CN_nD_E_SE_nSI, CN, nD, E, SE, nSI);
    and (CN_nD_E_nSE_SI, CN, nD, E, nSE, SI);
    and (CN_nD_E_nSE_nSI, CN, nD, E, nSE, nSI);
    and (nCN_D_E_SE_nSI, nCN, D, E, SE, nSI);
    and (nCN_D_E_nSE_SI, nCN, D, E, nSE, SI);
    and (nCN_D_E_nSE_nSI, nCN, D, E, nSE, nSI);
    and (nCN_D_nE_SE_nSI, nCN, D, nE, SE, nSI);
    and (nCN_D_nE_nSE_SI, nCN, D, nE, nSE, SI);
    and (nCN_D_nE_nSE_nSI, nCN, D, nE, nSE, nSI);
    and (nCN_nD_E_SE_nSI, nCN, nD, E, SE, nSI);
    and (nCN_nD_E_nSE_SI, nCN, nD, E, nSE, SI);
    and (nCN_nD_E_nSE_nSI, nCN, nD, E, nSE, nSI);
    and (nCN_nD_nE_SE_nSI, nCN, nD, nE, SE, nSI);
    and (nCN_nD_nE_nSE_SI, nCN, nD, nE, nSE, SI);
    and (nCN_nD_nE_nSE_nSI, nCN, nD, nE, nSE, nSI);
    and (CN_D_nE_SE_nSI, CN, D, nE, SE, nSI);
    and (CN_nD_nE_SE_nSI, CN, nD, nE, SE, nSI);
    and (D_E_nSE_SI, D, E, nSE, SI);
    and (D_E_nSE_nSI, D, E, nSE, nSI);
    and (D_nE_nSE_SI, D, nE, nSE, SI);
    and (D_nE_nSE_nSI, D, nE, nSE, nSI);
    and (nD_nE_nSE_SI, nD, nE, nSE, SI);
    and (nD_nE_nSE_nSI, nD, nE, nSE, nSI);
    and (CN_E_nSE_SI, CN, E, nSE, SI);
    and (CN_E_nSE_nSI, CN, E, nSE, nSI);
    and (CN_D_nSE_SI, CN, D, nSE, SI);
    and (CN_D_nSE_nSI, CN, D, nSE, nSI);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);
    and (CN_D_nE_SI, CN, D, nE, SI);
    and (CN_nD_nE_SI, CN, nD, nE, SI);
    and (CN_nD_E_SI, CN, nD, E, SI);
    and (nCN_D_E_SI, nCN, D, E, SI);
    and (nCN_D_nE_SI, nCN, D, nE, SI);
    and (nCN_nD_E_SI, nCN, nD, E, SI);
    and (nCN_nD_nE_SI, nCN, nD, nE, SI);
    and (CN_D_E_nSI, CN, D, E, nSI);
    and (CN_D_nE_nSI, CN, D, nE, nSI);
    and (CN_nD_nE_nSI, CN, nD, nE, nSI);
    and (CN_D_E_SE, CN, D, E, SE);
    and (CN_nD_E_SE, CN, nD, E, SE);
    and (nCN_D_E_SE, nCN, D, E, SE);
    and (nCN_D_nE_SE, nCN, D, nE, SE);
    and (nCN_nD_E_SE, nCN, nD, E, SE);
    and (nCN_nD_nE_SE, nCN, nD, nE, SE);
    and (CN_D_nE_SE, CN, D, nE, SE);
    and (CN_nD_nE_SE, CN, nD, nE, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    and  (D_check, E_d, CN_d, SE_int_not);
    and  (E_check, CN_d, SE_int_not);
    buf  (SI_check, SE_d);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    and  (D_check, E, CN, SE_int_not);
    and  (E_check, CN, SE_int_not);
    buf  (SI_check, SE);
  `endif
  buf  (CN_check, SE_int_not);
  or   (CP_check, D_check, E_check, CN_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && E && D) || (!(SE) && CN && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_E_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_E_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_E_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_E_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_E_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFKCNQD4 (SI, D, E, SE, CP, CN, Q);
    input SI, D, SE, CP, CN, E;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d, E_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        and (D2, CN_d, D1);
        tsmc_mux (D3, D2, SI_d, SE_d);
        tsmc_dff (Q_buf, D3, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        and (D2, CN, D1);
        tsmc_mux (D3, D2, SI, SE);
        tsmc_dff (Q_buf, D3, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_E_SE_SI_SDFCHK, CN_D_E_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_E_nSE_SI_SDFCHK, CN_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (CN_D_E_nSE_nSI_SDFCHK, CN_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_E_SE_SI_SDFCHK, CN_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nCN_D_E_SE_SI_SDFCHK, nCN_D_E_SE_SI, 1'b1);
    tsmc_xbuf (nCN_D_nE_SE_SI_SDFCHK, nCN_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_E_SE_SI_SDFCHK, nCN_nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SE_SI_SDFCHK, nCN_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_nE_SE_SI_SDFCHK, CN_D_nE_SE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nE_SE_SI_SDFCHK, CN_nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_E_SE_nSI_SDFCHK, CN_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_E_SE_nSI_SDFCHK, CN_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_E_nSE_SI_SDFCHK, CN_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_E_nSE_nSI_SDFCHK, CN_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_E_SE_nSI_SDFCHK, nCN_D_E_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_E_nSE_SI_SDFCHK, nCN_D_E_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_D_E_nSE_nSI_SDFCHK, nCN_D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_nE_SE_nSI_SDFCHK, nCN_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_nE_nSE_SI_SDFCHK, nCN_D_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_D_nE_nSE_nSI_SDFCHK, nCN_D_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_E_SE_nSI_SDFCHK, nCN_nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_E_nSE_SI_SDFCHK, nCN_nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_E_nSE_nSI_SDFCHK, nCN_nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SE_nSI_SDFCHK, nCN_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_nSE_SI_SDFCHK, nCN_nD_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_nSE_nSI_SDFCHK, nCN_nD_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_D_nE_SE_nSI_SDFCHK, CN_D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nE_SE_nSI_SDFCHK, CN_nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (D_E_nSE_SI_SDFCHK, D_E_nSE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_nSI_SDFCHK, D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nE_nSE_SI_SDFCHK, D_nE_nSE_SI, 1'b1);
    tsmc_xbuf (D_nE_nSE_nSI_SDFCHK, D_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_nSE_SI_SDFCHK, nD_nE_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nE_nSE_nSI_SDFCHK, nD_nE_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_E_nSE_SI_SDFCHK, CN_E_nSE_SI, 1'b1);
    tsmc_xbuf (CN_E_nSE_nSI_SDFCHK, CN_E_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SDFCHK, CN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SDFCHK, CN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_D_nE_SI_SDFCHK, CN_D_nE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nE_SI_SDFCHK, CN_nD_nE_SI, 1'b1);
    tsmc_xbuf (CN_nD_E_SI_SDFCHK, CN_nD_E_SI, 1'b1);
    tsmc_xbuf (nCN_D_E_SI_SDFCHK, nCN_D_E_SI, 1'b1);
    tsmc_xbuf (nCN_D_nE_SI_SDFCHK, nCN_D_nE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_E_SI_SDFCHK, nCN_nD_E_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SI_SDFCHK, nCN_nD_nE_SI, 1'b1);
    tsmc_xbuf (CN_D_E_nSI_SDFCHK, CN_D_E_nSI, 1'b1);
    tsmc_xbuf (CN_D_nE_nSI_SDFCHK, CN_D_nE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nE_nSI_SDFCHK, CN_nD_nE_nSI, 1'b1);
    tsmc_xbuf (CN_D_E_SE_SDFCHK, CN_D_E_SE, 1'b1);
    tsmc_xbuf (CN_nD_E_SE_SDFCHK, CN_nD_E_SE, 1'b1);
    tsmc_xbuf (nCN_D_E_SE_SDFCHK, nCN_D_E_SE, 1'b1);
    tsmc_xbuf (nCN_D_nE_SE_SDFCHK, nCN_D_nE_SE, 1'b1);
    tsmc_xbuf (nCN_nD_E_SE_SDFCHK, nCN_nD_E_SE, 1'b1);
    tsmc_xbuf (nCN_nD_nE_SE_SDFCHK, nCN_nD_nE_SE, 1'b1);
    tsmc_xbuf (CN_D_nE_SE_SDFCHK, CN_D_nE_SE, 1'b1);
    tsmc_xbuf (CN_nD_nE_SE_SDFCHK, CN_nD_nE_SE, 1'b1);
  `endif

    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    not (nE, E);
    and (CN_D_E_SE_SI, CN, D, E, SE, SI);
    and (CN_D_E_nSE_SI, CN, D, E, nSE, SI);
    and (CN_D_E_nSE_nSI, CN, D, E, nSE, nSI);
    and (CN_nD_E_SE_SI, CN, nD, E, SE, SI);
    and (nCN_D_E_SE_SI, nCN, D, E, SE, SI);
    and (nCN_D_nE_SE_SI, nCN, D, nE, SE, SI);
    and (nCN_nD_E_SE_SI, nCN, nD, E, SE, SI);
    and (nCN_nD_nE_SE_SI, nCN, nD, nE, SE, SI);
    and (CN_D_nE_SE_SI, CN, D, nE, SE, SI);
    and (CN_nD_nE_SE_SI, CN, nD, nE, SE, SI);
    and (CN_D_E_SE_nSI, CN, D, E, SE, nSI);
    and (CN_nD_E_SE_nSI, CN, nD, E, SE, nSI);
    and (CN_nD_E_nSE_SI, CN, nD, E, nSE, SI);
    and (CN_nD_E_nSE_nSI, CN, nD, E, nSE, nSI);
    and (nCN_D_E_SE_nSI, nCN, D, E, SE, nSI);
    and (nCN_D_E_nSE_SI, nCN, D, E, nSE, SI);
    and (nCN_D_E_nSE_nSI, nCN, D, E, nSE, nSI);
    and (nCN_D_nE_SE_nSI, nCN, D, nE, SE, nSI);
    and (nCN_D_nE_nSE_SI, nCN, D, nE, nSE, SI);
    and (nCN_D_nE_nSE_nSI, nCN, D, nE, nSE, nSI);
    and (nCN_nD_E_SE_nSI, nCN, nD, E, SE, nSI);
    and (nCN_nD_E_nSE_SI, nCN, nD, E, nSE, SI);
    and (nCN_nD_E_nSE_nSI, nCN, nD, E, nSE, nSI);
    and (nCN_nD_nE_SE_nSI, nCN, nD, nE, SE, nSI);
    and (nCN_nD_nE_nSE_SI, nCN, nD, nE, nSE, SI);
    and (nCN_nD_nE_nSE_nSI, nCN, nD, nE, nSE, nSI);
    and (CN_D_nE_SE_nSI, CN, D, nE, SE, nSI);
    and (CN_nD_nE_SE_nSI, CN, nD, nE, SE, nSI);
    and (D_E_nSE_SI, D, E, nSE, SI);
    and (D_E_nSE_nSI, D, E, nSE, nSI);
    and (D_nE_nSE_SI, D, nE, nSE, SI);
    and (D_nE_nSE_nSI, D, nE, nSE, nSI);
    and (nD_nE_nSE_SI, nD, nE, nSE, SI);
    and (nD_nE_nSE_nSI, nD, nE, nSE, nSI);
    and (CN_E_nSE_SI, CN, E, nSE, SI);
    and (CN_E_nSE_nSI, CN, E, nSE, nSI);
    and (CN_D_nSE_SI, CN, D, nSE, SI);
    and (CN_D_nSE_nSI, CN, D, nSE, nSI);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);
    and (CN_D_nE_SI, CN, D, nE, SI);
    and (CN_nD_nE_SI, CN, nD, nE, SI);
    and (CN_nD_E_SI, CN, nD, E, SI);
    and (nCN_D_E_SI, nCN, D, E, SI);
    and (nCN_D_nE_SI, nCN, D, nE, SI);
    and (nCN_nD_E_SI, nCN, nD, E, SI);
    and (nCN_nD_nE_SI, nCN, nD, nE, SI);
    and (CN_D_E_nSI, CN, D, E, nSI);
    and (CN_D_nE_nSI, CN, D, nE, nSI);
    and (CN_nD_nE_nSI, CN, nD, nE, nSI);
    and (CN_D_E_SE, CN, D, E, SE);
    and (CN_nD_E_SE, CN, nD, E, SE);
    and (nCN_D_E_SE, nCN, D, E, SE);
    and (nCN_D_nE_SE, nCN, D, nE, SE);
    and (nCN_nD_E_SE, nCN, nD, E, SE);
    and (nCN_nD_nE_SE, nCN, nD, nE, SE);
    and (CN_D_nE_SE, CN, D, nE, SE);
    and (CN_nD_nE_SE, CN, nD, nE, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    and  (D_check, E_d, CN_d, SE_int_not);
    and  (E_check, CN_d, SE_int_not);
    buf  (SI_check, SE_d);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    and  (D_check, E, CN, SE_int_not);
    and  (E_check, CN, SE_int_not);
    buf  (SI_check, SE);
  `endif
  buf  (CN_check, SE_int_not);
  or   (CP_check, D_check, E_check, CN_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && E && D) || (!(SE) && CN && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nE_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_E_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_E_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_E_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_E_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nE_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nE_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& CN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_E_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFQD0 (E, SE, CP, SI, D, Q);
    input E, SE, CP, SI, D;
    output Q;
    reg notifier;
    `ifdef NTC
        wire E_d, SE_d, CP_d, SI_d, D_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_E_SE_SI_SDFCHK, D_E_SE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_SI_SDFCHK, D_E_nSE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_nSI_SDFCHK, D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_E_SE_SI_SDFCHK, nD_E_SE_SI, 1'b1);
    tsmc_xbuf (D_nE_SE_SI_SDFCHK, D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SE_SI_SDFCHK, nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (D_E_SE_nSI_SDFCHK, D_E_SE_nSI, 1'b1);
    tsmc_xbuf (nD_E_SE_nSI_SDFCHK, nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (nD_E_nSE_SI_SDFCHK, nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (nD_E_nSE_nSI_SDFCHK, nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nE_SE_nSI_SDFCHK, D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_SE_nSI_SDFCHK, nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (E_nSE_SI_SDFCHK, E_nSE_SI, 1'b1);
    tsmc_xbuf (E_nSE_nSI_SDFCHK, E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nE_SI_SDFCHK, D_nE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SI_SDFCHK, nD_nE_SI, 1'b1);
    tsmc_xbuf (nD_E_SI_SDFCHK, nD_E_SI, 1'b1);
    tsmc_xbuf (D_E_nSI_SDFCHK, D_E_nSI, 1'b1);
    tsmc_xbuf (D_nE_nSI_SDFCHK, D_nE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_nSI_SDFCHK, nD_nE_nSI, 1'b1);
    tsmc_xbuf (D_E_SE_SDFCHK, D_E_SE, 1'b1);
    tsmc_xbuf (D_nE_SE_SDFCHK, D_nE_SE, 1'b1);
    tsmc_xbuf (nD_nE_SE_SDFCHK, nD_nE_SE, 1'b1);
    tsmc_xbuf (nD_E_SE_SDFCHK, nD_E_SE, 1'b1);
  `endif

    not (nE, E);
    not (nSE, SE);
    not (nSI, SI);
    not (nD, D);
    and (D_E_SE_SI, D, E, SE, SI);
    and (D_E_nSE_SI, D, E, nSE, SI);
    and (D_E_nSE_nSI, D, E, nSE, nSI);
    and (nD_E_SE_SI, nD, E, SE, SI);
    and (D_nE_SE_SI, D, nE, SE, SI);
    and (nD_nE_SE_SI, nD, nE, SE, SI);
    and (D_E_SE_nSI, D, E, SE, nSI);
    and (nD_E_SE_nSI, nD, E, SE, nSI);
    and (nD_E_nSE_SI, nD, E, nSE, SI);
    and (nD_E_nSE_nSI, nD, E, nSE, nSI);
    and (D_nE_SE_nSI, D, nE, SE, nSI);
    and (nD_nE_SE_nSI, nD, nE, SE, nSI);
    and (E_nSE_SI, E, nSE, SI);
    and (E_nSE_nSI, E, nSE, nSI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (D_nE_SI, D, nE, SI);
    and (nD_nE_SI, nD, nE, SI);
    and (nD_E_SI, nD, E, SI);
    and (D_E_nSI, D, E, nSI);
    and (D_nE_nSI, D, nE, nSI);
    and (nD_nE_nSI, nD, nE, nSI);
    and (D_E_SE, D, E, SE);
    and (D_nE_SE, D, nE, SE);
    and (nD_nE_SE, nD, nE, SE);
    and (nD_E_SE, nD, E, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFQD1 (E, SE, CP, SI, D, Q);
    input E, SE, CP, SI, D;
    output Q;
    reg notifier;
    `ifdef NTC
        wire E_d, SE_d, CP_d, SI_d, D_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_E_SE_SI_SDFCHK, D_E_SE_SI, 1'b1);
    tsmc_xbuf (D_nE_SE_SI_SDFCHK, D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nD_E_SE_SI_SDFCHK, nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SE_SI_SDFCHK, nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_SI_SDFCHK, D_E_nSE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_nSI_SDFCHK, D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_E_SE_nSI_SDFCHK, D_E_SE_nSI, 1'b1);
    tsmc_xbuf (D_nE_SE_nSI_SDFCHK, D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nD_E_SE_nSI_SDFCHK, nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_SE_nSI_SDFCHK, nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nD_E_nSE_SI_SDFCHK, nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (nD_E_nSE_nSI_SDFCHK, nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (E_nSE_SI_SDFCHK, E_nSE_SI, 1'b1);
    tsmc_xbuf (E_nSE_nSI_SDFCHK, E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nE_SI_SDFCHK, D_nE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SI_SDFCHK, nD_nE_SI, 1'b1);
    tsmc_xbuf (nD_E_SI_SDFCHK, nD_E_SI, 1'b1);
    tsmc_xbuf (D_E_nSI_SDFCHK, D_E_nSI, 1'b1);
    tsmc_xbuf (D_nE_nSI_SDFCHK, D_nE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_nSI_SDFCHK, nD_nE_nSI, 1'b1);
    tsmc_xbuf (D_E_SE_SDFCHK, D_E_SE, 1'b1);
    tsmc_xbuf (nD_E_SE_SDFCHK, nD_E_SE, 1'b1);
    tsmc_xbuf (D_nE_SE_SDFCHK, D_nE_SE, 1'b1);
    tsmc_xbuf (nD_nE_SE_SDFCHK, nD_nE_SE, 1'b1);
  `endif

    not (nE, E);
    not (nSE, SE);
    not (nSI, SI);
    not (nD, D);
    and (D_E_SE_SI, D, E, SE, SI);
    and (D_nE_SE_SI, D, nE, SE, SI);
    and (nD_E_SE_SI, nD, E, SE, SI);
    and (nD_nE_SE_SI, nD, nE, SE, SI);
    and (D_E_nSE_SI, D, E, nSE, SI);
    and (D_E_nSE_nSI, D, E, nSE, nSI);
    and (D_E_SE_nSI, D, E, SE, nSI);
    and (D_nE_SE_nSI, D, nE, SE, nSI);
    and (nD_E_SE_nSI, nD, E, SE, nSI);
    and (nD_nE_SE_nSI, nD, nE, SE, nSI);
    and (nD_E_nSE_SI, nD, E, nSE, SI);
    and (nD_E_nSE_nSI, nD, E, nSE, nSI);
    and (E_nSE_SI, E, nSE, SI);
    and (E_nSE_nSI, E, nSE, nSI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (D_nE_SI, D, nE, SI);
    and (nD_nE_SI, nD, nE, SI);
    and (nD_E_SI, nD, E, SI);
    and (D_E_nSI, D, E, nSI);
    and (D_nE_nSI, D, nE, nSI);
    and (nD_nE_nSI, nD, nE, nSI);
    and (D_E_SE, D, E, SE);
    and (nD_E_SE, nD, E, SE);
    and (D_nE_SE, D, nE, SE);
    and (nD_nE_SE, nD, nE, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFQD2 (E, SE, CP, SI, D, Q);
    input E, SE, CP, SI, D;
    output Q;
    reg notifier;
    `ifdef NTC
        wire E_d, SE_d, CP_d, SI_d, D_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_E_SE_SI_SDFCHK, D_E_SE_SI, 1'b1);
    tsmc_xbuf (D_nE_SE_SI_SDFCHK, D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nD_E_SE_SI_SDFCHK, nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SE_SI_SDFCHK, nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_SI_SDFCHK, D_E_nSE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_nSI_SDFCHK, D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_E_SE_nSI_SDFCHK, D_E_SE_nSI, 1'b1);
    tsmc_xbuf (D_nE_SE_nSI_SDFCHK, D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nD_E_SE_nSI_SDFCHK, nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_SE_nSI_SDFCHK, nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nD_E_nSE_SI_SDFCHK, nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (nD_E_nSE_nSI_SDFCHK, nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (E_nSE_SI_SDFCHK, E_nSE_SI, 1'b1);
    tsmc_xbuf (E_nSE_nSI_SDFCHK, E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nE_SI_SDFCHK, D_nE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SI_SDFCHK, nD_nE_SI, 1'b1);
    tsmc_xbuf (nD_E_SI_SDFCHK, nD_E_SI, 1'b1);
    tsmc_xbuf (D_E_nSI_SDFCHK, D_E_nSI, 1'b1);
    tsmc_xbuf (D_nE_nSI_SDFCHK, D_nE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_nSI_SDFCHK, nD_nE_nSI, 1'b1);
    tsmc_xbuf (D_E_SE_SDFCHK, D_E_SE, 1'b1);
    tsmc_xbuf (nD_E_SE_SDFCHK, nD_E_SE, 1'b1);
    tsmc_xbuf (D_nE_SE_SDFCHK, D_nE_SE, 1'b1);
    tsmc_xbuf (nD_nE_SE_SDFCHK, nD_nE_SE, 1'b1);
  `endif

    not (nE, E);
    not (nSE, SE);
    not (nSI, SI);
    not (nD, D);
    and (D_E_SE_SI, D, E, SE, SI);
    and (D_nE_SE_SI, D, nE, SE, SI);
    and (nD_E_SE_SI, nD, E, SE, SI);
    and (nD_nE_SE_SI, nD, nE, SE, SI);
    and (D_E_nSE_SI, D, E, nSE, SI);
    and (D_E_nSE_nSI, D, E, nSE, nSI);
    and (D_E_SE_nSI, D, E, SE, nSI);
    and (D_nE_SE_nSI, D, nE, SE, nSI);
    and (nD_E_SE_nSI, nD, E, SE, nSI);
    and (nD_nE_SE_nSI, nD, nE, SE, nSI);
    and (nD_E_nSE_SI, nD, E, nSE, SI);
    and (nD_E_nSE_nSI, nD, E, nSE, nSI);
    and (E_nSE_SI, E, nSE, SI);
    and (E_nSE_nSI, E, nSE, nSI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (D_nE_SI, D, nE, SI);
    and (nD_nE_SI, nD, nE, SI);
    and (nD_E_SI, nD, E, SI);
    and (D_E_nSI, D, E, nSI);
    and (D_nE_nSI, D, nE, nSI);
    and (nD_nE_nSI, nD, nE, nSI);
    and (D_E_SE, D, E, SE);
    and (nD_E_SE, nD, E, SE);
    and (D_nE_SE, D, nE, SE);
    and (nD_nE_SE, nD, nE, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFQD4 (E, SE, CP, SI, D, Q);
    input E, SE, CP, SI, D;
    output Q;
    reg notifier;
    `ifdef NTC
        wire E_d, SE_d, CP_d, SI_d, D_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_E_SE_SI_SDFCHK, D_E_SE_SI, 1'b1);
    tsmc_xbuf (D_nE_SE_SI_SDFCHK, D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nD_E_SE_SI_SDFCHK, nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SE_SI_SDFCHK, nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_SI_SDFCHK, D_E_nSE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_nSI_SDFCHK, D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_E_SE_nSI_SDFCHK, D_E_SE_nSI, 1'b1);
    tsmc_xbuf (D_nE_SE_nSI_SDFCHK, D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nD_E_SE_nSI_SDFCHK, nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_SE_nSI_SDFCHK, nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nD_E_nSE_SI_SDFCHK, nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (nD_E_nSE_nSI_SDFCHK, nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (E_nSE_SI_SDFCHK, E_nSE_SI, 1'b1);
    tsmc_xbuf (E_nSE_nSI_SDFCHK, E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nE_SI_SDFCHK, D_nE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SI_SDFCHK, nD_nE_SI, 1'b1);
    tsmc_xbuf (nD_E_SI_SDFCHK, nD_E_SI, 1'b1);
    tsmc_xbuf (D_E_nSI_SDFCHK, D_E_nSI, 1'b1);
    tsmc_xbuf (D_nE_nSI_SDFCHK, D_nE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_nSI_SDFCHK, nD_nE_nSI, 1'b1);
    tsmc_xbuf (D_E_SE_SDFCHK, D_E_SE, 1'b1);
    tsmc_xbuf (nD_E_SE_SDFCHK, nD_E_SE, 1'b1);
    tsmc_xbuf (D_nE_SE_SDFCHK, D_nE_SE, 1'b1);
    tsmc_xbuf (nD_nE_SE_SDFCHK, nD_nE_SE, 1'b1);
  `endif

    not (nE, E);
    not (nSE, SE);
    not (nSI, SI);
    not (nD, D);
    and (D_E_SE_SI, D, E, SE, SI);
    and (D_nE_SE_SI, D, nE, SE, SI);
    and (nD_E_SE_SI, nD, E, SE, SI);
    and (nD_nE_SE_SI, nD, nE, SE, SI);
    and (D_E_nSE_SI, D, E, nSE, SI);
    and (D_E_nSE_nSI, D, E, nSE, nSI);
    and (D_E_SE_nSI, D, E, SE, nSI);
    and (D_nE_SE_nSI, D, nE, SE, nSI);
    and (nD_E_SE_nSI, nD, E, SE, nSI);
    and (nD_nE_SE_nSI, nD, nE, SE, nSI);
    and (nD_E_nSE_SI, nD, E, nSE, SI);
    and (nD_E_nSE_nSI, nD, E, nSE, nSI);
    and (E_nSE_SI, E, nSE, SI);
    and (E_nSE_nSI, E, nSE, nSI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (D_nE_SI, D, nE, SI);
    and (nD_nE_SI, nD, nE, SI);
    and (nD_E_SI, nD, E, SI);
    and (D_E_nSI, D, E, nSI);
    and (D_nE_nSI, D, nE, nSI);
    and (nD_nE_nSI, nD, nE, nSI);
    and (D_E_SE, D, E, SE);
    and (nD_E_SE, nD, E, SE);
    and (D_nE_SE, D, nE, SE);
    and (nD_nE_SE, nD, nE, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFQND0 (E, SE, CP, SI, D, QN);
    input E, SE, CP, SI, D;
    output QN;
    reg notifier;
    `ifdef NTC
        wire E_d, SE_d, CP_d, SI_d, D_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_E_SE_nSI_SDFCHK, D_E_SE_nSI, 1'b1);
    tsmc_xbuf (nD_E_SE_nSI_SDFCHK, nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (nD_E_nSE_SI_SDFCHK, nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (nD_E_nSE_nSI_SDFCHK, nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nE_SE_nSI_SDFCHK, D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_SE_nSI_SDFCHK, nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (D_E_SE_SI_SDFCHK, D_E_SE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_SI_SDFCHK, D_E_nSE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_nSI_SDFCHK, D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_E_SE_SI_SDFCHK, nD_E_SE_SI, 1'b1);
    tsmc_xbuf (D_nE_SE_SI_SDFCHK, D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SE_SI_SDFCHK, nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (E_nSE_SI_SDFCHK, E_nSE_SI, 1'b1);
    tsmc_xbuf (E_nSE_nSI_SDFCHK, E_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (D_E_nSI_SDFCHK, D_E_nSI, 1'b1);
    tsmc_xbuf (D_nE_nSI_SDFCHK, D_nE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_nSI_SDFCHK, nD_nE_nSI, 1'b1);
    tsmc_xbuf (D_nE_SI_SDFCHK, D_nE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SI_SDFCHK, nD_nE_SI, 1'b1);
    tsmc_xbuf (nD_E_SI_SDFCHK, nD_E_SI, 1'b1);
    tsmc_xbuf (D_E_SE_SDFCHK, D_E_SE, 1'b1);
    tsmc_xbuf (D_nE_SE_SDFCHK, D_nE_SE, 1'b1);
    tsmc_xbuf (nD_nE_SE_SDFCHK, nD_nE_SE, 1'b1);
    tsmc_xbuf (nD_E_SE_SDFCHK, nD_E_SE, 1'b1);
  `endif

    not (nE, E);
    not (nSE, SE);
    not (nSI, SI);
    not (nD, D);
    and (D_E_SE_nSI, D, E, SE, nSI);
    and (nD_E_SE_nSI, nD, E, SE, nSI);
    and (nD_E_nSE_SI, nD, E, nSE, SI);
    and (nD_E_nSE_nSI, nD, E, nSE, nSI);
    and (D_nE_SE_nSI, D, nE, SE, nSI);
    and (nD_nE_SE_nSI, nD, nE, SE, nSI);
    and (D_E_SE_SI, D, E, SE, SI);
    and (D_E_nSE_SI, D, E, nSE, SI);
    and (D_E_nSE_nSI, D, E, nSE, nSI);
    and (nD_E_SE_SI, nD, E, SE, SI);
    and (D_nE_SE_SI, D, nE, SE, SI);
    and (nD_nE_SE_SI, nD, nE, SE, SI);
    and (E_nSE_SI, E, nSE, SI);
    and (E_nSE_nSI, E, nSE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (D_E_nSI, D, E, nSI);
    and (D_nE_nSI, D, nE, nSI);
    and (nD_nE_nSI, nD, nE, nSI);
    and (D_nE_SI, D, nE, SI);
    and (nD_nE_SI, nD, nE, SI);
    and (nD_E_SI, nD, E, SI);
    and (D_E_SE, D, E, SE);
    and (D_nE_SE, D, nE, SE);
    and (nD_nE_SE, nD, nE, SE);
    and (nD_E_SE, nD, E, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (QN-:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFQND1 (E, SE, CP, SI, D, QN);
    input E, SE, CP, SI, D;
    output QN;
    reg notifier;
    `ifdef NTC
        wire E_d, SE_d, CP_d, SI_d, D_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_E_SE_nSI_SDFCHK, D_E_SE_nSI, 1'b1);
    tsmc_xbuf (D_nE_SE_nSI_SDFCHK, D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nD_E_SE_nSI_SDFCHK, nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_SE_nSI_SDFCHK, nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nD_E_nSE_SI_SDFCHK, nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (nD_E_nSE_nSI_SDFCHK, nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_E_SE_SI_SDFCHK, D_E_SE_SI, 1'b1);
    tsmc_xbuf (D_nE_SE_SI_SDFCHK, D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nD_E_SE_SI_SDFCHK, nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SE_SI_SDFCHK, nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_SI_SDFCHK, D_E_nSE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_nSI_SDFCHK, D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (E_nSE_SI_SDFCHK, E_nSE_SI, 1'b1);
    tsmc_xbuf (E_nSE_nSI_SDFCHK, E_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (D_E_nSI_SDFCHK, D_E_nSI, 1'b1);
    tsmc_xbuf (D_nE_nSI_SDFCHK, D_nE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_nSI_SDFCHK, nD_nE_nSI, 1'b1);
    tsmc_xbuf (D_nE_SI_SDFCHK, D_nE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SI_SDFCHK, nD_nE_SI, 1'b1);
    tsmc_xbuf (nD_E_SI_SDFCHK, nD_E_SI, 1'b1);
    tsmc_xbuf (D_E_SE_SDFCHK, D_E_SE, 1'b1);
    tsmc_xbuf (nD_E_SE_SDFCHK, nD_E_SE, 1'b1);
    tsmc_xbuf (D_nE_SE_SDFCHK, D_nE_SE, 1'b1);
    tsmc_xbuf (nD_nE_SE_SDFCHK, nD_nE_SE, 1'b1);
  `endif

    not (nE, E);
    not (nSE, SE);
    not (nSI, SI);
    not (nD, D);
    and (D_E_SE_nSI, D, E, SE, nSI);
    and (D_nE_SE_nSI, D, nE, SE, nSI);
    and (nD_E_SE_nSI, nD, E, SE, nSI);
    and (nD_nE_SE_nSI, nD, nE, SE, nSI);
    and (nD_E_nSE_SI, nD, E, nSE, SI);
    and (nD_E_nSE_nSI, nD, E, nSE, nSI);
    and (D_E_SE_SI, D, E, SE, SI);
    and (D_nE_SE_SI, D, nE, SE, SI);
    and (nD_E_SE_SI, nD, E, SE, SI);
    and (nD_nE_SE_SI, nD, nE, SE, SI);
    and (D_E_nSE_SI, D, E, nSE, SI);
    and (D_E_nSE_nSI, D, E, nSE, nSI);
    and (E_nSE_SI, E, nSE, SI);
    and (E_nSE_nSI, E, nSE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (D_E_nSI, D, E, nSI);
    and (D_nE_nSI, D, nE, nSI);
    and (nD_nE_nSI, nD, nE, nSI);
    and (D_nE_SI, D, nE, SI);
    and (nD_nE_SI, nD, nE, SI);
    and (nD_E_SI, nD, E, SI);
    and (D_E_SE, D, E, SE);
    and (nD_E_SE, nD, E, SE);
    and (D_nE_SE, D, nE, SE);
    and (nD_nE_SE, nD, nE, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (QN-:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFQND2 (E, SE, CP, SI, D, QN);
    input E, SE, CP, SI, D;
    output QN;
    reg notifier;
    `ifdef NTC
        wire E_d, SE_d, CP_d, SI_d, D_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_E_SE_nSI_SDFCHK, D_E_SE_nSI, 1'b1);
    tsmc_xbuf (D_nE_SE_nSI_SDFCHK, D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nD_E_SE_nSI_SDFCHK, nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_SE_nSI_SDFCHK, nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nD_E_nSE_SI_SDFCHK, nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (nD_E_nSE_nSI_SDFCHK, nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_E_SE_SI_SDFCHK, D_E_SE_SI, 1'b1);
    tsmc_xbuf (D_nE_SE_SI_SDFCHK, D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nD_E_SE_SI_SDFCHK, nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SE_SI_SDFCHK, nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_SI_SDFCHK, D_E_nSE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_nSI_SDFCHK, D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (E_nSE_SI_SDFCHK, E_nSE_SI, 1'b1);
    tsmc_xbuf (E_nSE_nSI_SDFCHK, E_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (D_E_nSI_SDFCHK, D_E_nSI, 1'b1);
    tsmc_xbuf (D_nE_nSI_SDFCHK, D_nE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_nSI_SDFCHK, nD_nE_nSI, 1'b1);
    tsmc_xbuf (D_nE_SI_SDFCHK, D_nE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SI_SDFCHK, nD_nE_SI, 1'b1);
    tsmc_xbuf (nD_E_SI_SDFCHK, nD_E_SI, 1'b1);
    tsmc_xbuf (D_E_SE_SDFCHK, D_E_SE, 1'b1);
    tsmc_xbuf (nD_E_SE_SDFCHK, nD_E_SE, 1'b1);
    tsmc_xbuf (D_nE_SE_SDFCHK, D_nE_SE, 1'b1);
    tsmc_xbuf (nD_nE_SE_SDFCHK, nD_nE_SE, 1'b1);
  `endif

    not (nE, E);
    not (nSE, SE);
    not (nSI, SI);
    not (nD, D);
    and (D_E_SE_nSI, D, E, SE, nSI);
    and (D_nE_SE_nSI, D, nE, SE, nSI);
    and (nD_E_SE_nSI, nD, E, SE, nSI);
    and (nD_nE_SE_nSI, nD, nE, SE, nSI);
    and (nD_E_nSE_SI, nD, E, nSE, SI);
    and (nD_E_nSE_nSI, nD, E, nSE, nSI);
    and (D_E_SE_SI, D, E, SE, SI);
    and (D_nE_SE_SI, D, nE, SE, SI);
    and (nD_E_SE_SI, nD, E, SE, SI);
    and (nD_nE_SE_SI, nD, nE, SE, SI);
    and (D_E_nSE_SI, D, E, nSE, SI);
    and (D_E_nSE_nSI, D, E, nSE, nSI);
    and (E_nSE_SI, E, nSE, SI);
    and (E_nSE_nSI, E, nSE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (D_E_nSI, D, E, nSI);
    and (D_nE_nSI, D, nE, nSI);
    and (nD_nE_nSI, nD, nE, nSI);
    and (D_nE_SI, D, nE, SI);
    and (nD_nE_SI, nD, nE, SI);
    and (nD_E_SI, nD, E, SI);
    and (D_E_SE, D, E, SE);
    and (nD_E_SE, nD, E, SE);
    and (D_nE_SE, D, nE, SE);
    and (nD_nE_SE, nD, nE, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (QN-:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFQND4 (E, SE, CP, SI, D, QN);
    input E, SE, CP, SI, D;
    output QN;
    reg notifier;
    `ifdef NTC
        wire E_d, SE_d, CP_d, SI_d, D_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D_d, E_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D1, Q_buf, D, E);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_E_SE_nSI_SDFCHK, D_E_SE_nSI, 1'b1);
    tsmc_xbuf (D_nE_SE_nSI_SDFCHK, D_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nD_E_SE_nSI_SDFCHK, nD_E_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_SE_nSI_SDFCHK, nD_nE_SE_nSI, 1'b1);
    tsmc_xbuf (nD_E_nSE_SI_SDFCHK, nD_E_nSE_SI, 1'b1);
    tsmc_xbuf (nD_E_nSE_nSI_SDFCHK, nD_E_nSE_nSI, 1'b1);
    tsmc_xbuf (D_E_SE_SI_SDFCHK, D_E_SE_SI, 1'b1);
    tsmc_xbuf (D_nE_SE_SI_SDFCHK, D_nE_SE_SI, 1'b1);
    tsmc_xbuf (nD_E_SE_SI_SDFCHK, nD_E_SE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SE_SI_SDFCHK, nD_nE_SE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_SI_SDFCHK, D_E_nSE_SI, 1'b1);
    tsmc_xbuf (D_E_nSE_nSI_SDFCHK, D_E_nSE_nSI, 1'b1);
    tsmc_xbuf (E_nSE_SI_SDFCHK, E_nSE_SI, 1'b1);
    tsmc_xbuf (E_nSE_nSI_SDFCHK, E_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (D_E_nSI_SDFCHK, D_E_nSI, 1'b1);
    tsmc_xbuf (D_nE_nSI_SDFCHK, D_nE_nSI, 1'b1);
    tsmc_xbuf (nD_nE_nSI_SDFCHK, nD_nE_nSI, 1'b1);
    tsmc_xbuf (D_nE_SI_SDFCHK, D_nE_SI, 1'b1);
    tsmc_xbuf (nD_nE_SI_SDFCHK, nD_nE_SI, 1'b1);
    tsmc_xbuf (nD_E_SI_SDFCHK, nD_E_SI, 1'b1);
    tsmc_xbuf (D_E_SE_SDFCHK, D_E_SE, 1'b1);
    tsmc_xbuf (nD_E_SE_SDFCHK, nD_E_SE, 1'b1);
    tsmc_xbuf (D_nE_SE_SDFCHK, D_nE_SE, 1'b1);
    tsmc_xbuf (nD_nE_SE_SDFCHK, nD_nE_SE, 1'b1);
  `endif

    not (nE, E);
    not (nSE, SE);
    not (nSI, SI);
    not (nD, D);
    and (D_E_SE_nSI, D, E, SE, nSI);
    and (D_nE_SE_nSI, D, nE, SE, nSI);
    and (nD_E_SE_nSI, nD, E, SE, nSI);
    and (nD_nE_SE_nSI, nD, nE, SE, nSI);
    and (nD_E_nSE_SI, nD, E, nSE, SI);
    and (nD_E_nSE_nSI, nD, E, nSE, nSI);
    and (D_E_SE_SI, D, E, SE, SI);
    and (D_nE_SE_SI, D, nE, SE, SI);
    and (nD_E_SE_SI, nD, E, SE, SI);
    and (nD_nE_SE_SI, nD, nE, SE, SI);
    and (D_E_nSE_SI, D, E, nSE, SI);
    and (D_E_nSE_nSI, D, E, nSE, nSI);
    and (E_nSE_SI, E, nSE, SI);
    and (E_nSE_nSI, E, nSE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (D_E_nSI, D, E, nSI);
    and (D_nE_nSI, D, nE, nSI);
    and (nD_nE_nSI, nD, nE, nSI);
    and (D_nE_SI, D, nE, SI);
    and (nD_nE_SI, nD, nE, SI);
    and (nD_E_SI, nD, E, SI);
    and (D_E_SE, D, E, SE);
    and (nD_E_SE, nD, E, SE);
    and (D_nE_SE, D, nE, SE);
    and (nD_nE_SE, nD, nE, SE);

  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (QN-:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nE_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_E_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nE_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_E_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& E_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_E_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nE_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module TIEH (Z);
    output Z;
    buf (Z, 1'b1);

endmodule
`endcelldefine

`celldefine
module TIEL (ZN);
    output ZN;
    buf (ZN, 1'b0);

endmodule
`endcelldefine

`celldefine
module XNR2D0 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    xor (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    if (A2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0)
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR2D1 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    xor (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    if (A2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0)
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR2D2 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    xor (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    if (A2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0)
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR2D4 (A1, A2, ZN);
    input A1, A2;
    output ZN;
    xor (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    if (A2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0)
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR3D0 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    xor (I0_out, A1, A2);
    xor (I1_out, I0_out, A3);
    not (ZN, I1_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR3D1 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    xor (I0_out, A1, A2);
    xor (I1_out, I0_out, A3);
    not (ZN, I1_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR3D2 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    xor (I0_out, A1, A2);
    xor (I1_out, I0_out, A3);
    not (ZN, I1_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR3D4 (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    xor (I0_out, A1, A2);
    xor (I1_out, I0_out, A3);
    not (ZN, I1_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR4D0 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    xor (I0_out, A1, A2);
    xor (I1_out, I0_out, A3);
    xor (I2_out, I1_out, A4);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR4D1 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    xor (I0_out, A1, A2);
    xor (I1_out, I0_out, A3);
    xor (I2_out, I1_out, A4);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR4D2 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    xor (I0_out, A1, A2);
    xor (I1_out, I0_out, A3);
    xor (I2_out, I1_out, A4);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR4D4 (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    xor (I0_out, A1, A2);
    xor (I1_out, I0_out, A3);
    xor (I2_out, I1_out, A4);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR2D0 (A1, A2, Z);
    input A1, A2;
    output Z;
    xor (Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR2D1 (A1, A2, Z);
    input A1, A2;
    output Z;
    xor (Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR2D2 (A1, A2, Z);
    input A1, A2;
    output Z;
    xor (Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR2D4 (A1, A2, Z);
    input A1, A2;
    output Z;
    xor (Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR3D0 (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    xor (I0_out, A1, A2);
    xor (Z, I0_out, A3);

  specify
    if (A2 == 1'b1 && A3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR3D1 (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    xor (I0_out, A1, A2);
    xor (Z, I0_out, A3);

  specify
    if (A2 == 1'b1 && A3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR3D2 (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    xor (I0_out, A1, A2);
    xor (Z, I0_out, A3);

  specify
    if (A2 == 1'b1 && A3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR3D4 (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    xor (I0_out, A1, A2);
    xor (Z, I0_out, A3);

  specify
    if (A2 == 1'b1 && A3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR4D0 (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    xor (I0_out, A1, A2);
    xor (I1_out, I0_out, A3);
    xor (Z, I1_out, A4);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR4D1 (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    xor (I0_out, A1, A2);
    xor (I1_out, I0_out, A3);
    xor (Z, I1_out, A4);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR4D2 (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    xor (I0_out, A1, A2);
    xor (I1_out, I0_out, A3);
    xor (Z, I1_out, A4);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR4D4 (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    xor (I0_out, A1, A2);
    xor (I1_out, I0_out, A3);
    xor (Z, I1_out, A4);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

primitive tsmc_mux (q, d0, d1, s);
   output q;
   input s, d0, d1;

   table
   // d0  d1  s   : q 
      0   ?   0   : 0 ;
      1   ?   0   : 1 ;
      ?   0   1   : 0 ;
      ?   1   1   : 1 ;
      0   0   x   : 0 ;
      1   1   x   : 1 ;
   endtable
endprimitive
primitive tsmc_dla (q, d, e, cdn, sdn, notifier);
   output q;
   reg q;
   input d, e, cdn, sdn, notifier;
   table
   1  1   1   ?   ?   : ?  :  1  ; // Latch 1
   0  1   ?   1   ?   : ?  :  0  ; // Latch 0
   0 (10) 1   1   ?   : ?  :  0  ; // Latch 0 after falling edge
   1 (10) 1   1   ?   : ?  :  1  ; // Latch 1 after falling edge
   *  0   ?   ?   ?   : ?  :  -  ; // no changes
   ?  ?   ?   0   ?   : ?  :  1  ; // preset to 1
   ?  0   1   *   ?   : 1  :  1  ;
   1  ?   1   *   ?   : 1  :  1  ;
   1  *   1   ?   ?   : 1  :  1  ;
   ?  ?   0   1   ?   : ?  :  0  ; // reset to 0
   ?  0   *   1   ?   : 0  :  0  ;
   0  ?   *   1   ?   : 0  :  0  ;
   0  *   ?   1   ?   : 0  :  0  ;
   ?  ?   ?   ?   *   : ?  :  x  ; // toggle notifier
   endtable
endprimitive
primitive tsmc_xbuf (o, i, dummy);
   output o;     
   input i, dummy;
   table         
   // i dummy : o
      0   1   : 0 ;
      1   1   : 1 ;
      x   1   : 1 ;
   endtable      
endprimitive 
primitive tsmc_dff (q, d, cp, cdn, sdn, notifier);
   output q;
   input d, cp, cdn, sdn, notifier;
   reg q;
   table
      ?   ?   0   ?   ? : ? : 0 ; // CDN dominate SDN
      ?   ?   1   0   ? : ? : 1 ; // SDN is set   
      ?   ?   1   x   ? : 0 : x ; // SDN affect Q
      ?   ?   1   x   ? : 1 : 1 ; // Q=1,preset=X
      ?   ?   x   1   ? : 0 : 0 ; // Q=0,clear=X
      0 (01)  ?   1   ? : ? : 0 ; // Latch 0
      0 (0x)  1   1   ? : ? : x ; // Weak clock
      0   0   ?   1   ? : 0 : 0 ; // Keep 0 (D==Q)
      1 (01)  1   ?   ? : ? : 1 ; // Latch 1   
      1 (0x)  1   ?   ? : ? : x ; // Weak clock
      1   0   1   ?   ? : 1 : 1 ; // Keep 1 (D==Q)
      ? (1?)  1   1   ? : ? : - ; // ignore negative edge of clock
      ?   0   1   1   ? : ? : - ; // ignore low-level clock
      ?   ? (?1)  1   ? : ? : - ; // ignore positive edge of CDN
      ?   ?   1 (?1)  ? : ? : - ; // ignore posative edge of SDN
      *   ?   1   1   ? : ? : - ; // ignore data change on steady clock
      ?   ?   ?   ?   * : ? : x ; // timing check violation
   endtable
endprimitive
